`default_nettype none

module tt_um_adpll (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
  //assign uo_out  = 0;  // Example: ou_out is the sum of ui_in and uio_in
  assign uio_out = 0;
  assign uio_oe  = 0;
  // List all unused inputs to prevent warnings
	wire _unused = &{ena,uio_in,1'b0};
   adpll adp(
    .vco_clk(clk),
    .clk2_5k(ui_in[0]),
    .tdc_reset(rst_n),   
    .out(uo_out[5]),
    .vco_in(uo_out[3:0]),
    .desired_out(uo_out[4])
    );
  endmodule
module adpll(vco_clk, clk2_5k, tdc_reset, out, vco_in,desired_out);
	input tdc_reset;
	input vco_clk,clk2_5k;// clk2_5k;
	output out;// clk2_5k;
	output desired_out;
	output [3:0] vco_in;
	wire [15:0] s;
	wire [15:0] t;
	wire freq_div_out;
	wire [3:0] encoder_out;
	
	// FLASH TDC with resolution = 24 us 
	tdc_in m1(tdc_reset, vco_clk, freq_div_out, s);
	tdc_ref m2(clk2_5k, s, t);
	
	// Produces VCO_IN based on the digital code obtained from TDC
	encoder m3(t, encoder_out);
	dlf m4(encoder_out, vco_in, clk2_5k);
	
	// Works on 50 MHz and provides the 16 frequencies from 2 KHz to 17 KHz
	vco m5(vco_clk, vco_in, out, desired_out);
	
	// Divide by 4 frequency divider
	freq_div m6(out, freq_div_out); 
endmodule

module tdc_in(tdc_reset, vco_clk, clk, out);
	input tdc_reset, vco_clk, clk;
	output reg [15:0] out=0;
//	integer i = 0; 
	wire en = 1;
	wire [11:0] sin_out, cos_out, squ_out;
	wire wave_out;
	wire ref24;
	

	waveform_gen dut (
    .clk(vco_clk),
    .reset(tdc_reset),
    .en(en),
    .phase_inc(32'h00038FCE2),//369D03), // to generate 24us signal which is the resolution of our TDC
    .sin_out(sin_out),
	 .cos_out(cos_out),
    .squ_out(squ_out),
	 .vco_out(ref24),
	 .desired_freq_sig(wave_out)
);
	
	always@(posedge ref24)
	begin
		out[0] <= clk;
		out[1] <= out[0];
		out[2] <= out[1];
		out[3] <= out[2];
		out[4] <= out[3];
		out[5] <= out[4];
		out[6] <= out[5];
		out[7] <= out[6];
		out[8] <= out[7];
		out[9] <= out[8];
		out[10] <= out[9];
		out[11] <= out[10];
		out[12] <= out[11];
		out[13] <= out[12];
		out[14] <= out[13];
		out[15] <= out[14];
	end
//	
endmodule

module tdc_ref(clk, in, out);
	input clk;
	input [15:0] in;
	output reg [15:0] out=0;
	integer i = 0;
	always@(posedge clk)
	begin
		for(i=0; i<16; i = i + 1)
		begin
			out[i] <= in[i];
		end
	end
endmodule

module encoder (in, out);
	input [15:0] in;
	output reg [3:0] out = 0;    
	always@(*)
	begin  
		if((16'hffff & in) == 16'hffff) out = 4'b0111;
		else if((16'h7fff & in) == 16'h7fff) out = 4'b0111;
		else if((16'h3fff & in) == 16'h3fff) out = 4'b0110;
		else if((16'h1fff & in) == 16'h1fff) out = 4'b0101;
		else if((16'h0fff & in) == 16'h0fff) out = 4'b0100;
		else if((16'h07ff & in) == 16'h07ff) out = 4'b0011;
		else if((16'h03ff & in) == 16'h03ff) out = 4'b0010;
		else if((16'h01ff & in) == 16'h01ff) out = 4'b0001;
		else if((16'h00ff & in) == 16'h00ff) out = 4'b1111;
		else if((16'h007f & in) == 16'h007f) out = 4'b1110;
		else if((16'h003f & in) == 16'h003f) out = 4'b1101;
		else if((16'h001f & in) == 16'h001f) out = 4'b1100;
		else if((16'h000f & in) == 16'h000f) out = 4'b1011;
		else if((16'h0007 & in) == 16'h0007) out = 4'b1010;
		else if((16'h0003 & in) == 16'h0003) out = 4'b1001;
		else if((16'h0001 & in) == 16'h0001) out = 4'b1000;
		else out = 4'b0000;
	end 
endmodule

module dlf (in, out, clk);
	input clk;
	input signed [3:0] in;
	output [3:0] out;
//	wire signed [3:0] acc;   ///original filter
//	reg signed [3:0] latch = 0; 
//	parameter a = 1;// b = 1;
//	assign acc = latch + (in >>> 2); //in/4
//	//assign out = acc + (in * a);
//	assign out = acc + in; //same as a=1 ?
//	always@(posedge clk)
//	begin
//		latch <= acc;
//	end


reg signed [3:0] latch1 = 0; // moving summation filter
reg signed [3:0] latch2 = 0;
reg signed [3:0] latch3 = 0;
wire signed [3:0] acc;

	always@(posedge clk)
	begin
		latch1 <= in;
	end
	
	always@(posedge clk)
	begin
		latch2 <= latch1;
	end	
	
	always@(posedge clk)
	begin
		latch3 <= latch2;
	end
	
	assign acc = latch1 + latch2 + latch3 +in;
	
	assign out= (acc>>0);

//	reg signed [3:0] latch1 = 0; // IIR filter
//reg signed [3:0] latch2 = 0;
//wire signed [3:0] acc;
//wire signed [3:0] shifter;
//	
//	always@(posedge clk)
//	begin
//		latch1 <= in;
//	end
//	
//	assign acc = latch1 + in;
//	
//	always@(posedge clk)
//	begin
//		latch2 <= out;
//	end	
//	
//	assign shifter=(latch2>>2);
//	
//	assign out=(shifter*4'd3)+acc;
endmodule 

module vco (vco_clk, in, out, desired_out);
   input vco_clk;
//	input reset;
	input [3:0] in;
	output wire out;
	output wire desired_out;
	
	reg [31:0] phase_inc;
	wire en=1;
	reg reset;
	reg [3:0]in_reg;
	wire got_it;
	wire [11:0] sin_out;
	wire [11:0] cos_out;
	wire [11:0] squ_out;
waveform_gen dut (
    .clk(vco_clk),
    .reset(reset),
    .en(en),
    .phase_inc(phase_inc),
    .sin_out(sin_out),
	 .cos_out(cos_out),
    .squ_out(squ_out),
	 .vco_out(out),
	 .desired_freq_sig(desired_out)
);

always@(posedge vco_clk)
	begin
		in_reg <= in;
		if((in_reg == in))
			reset <= 1;
		else
			reset <= 0;
	end

always@(*)
	begin
	//with VCO CLOCK = 50 MHz

		case (in)
			4'h0 :
			begin
				phase_inc = 32'h00029F16;//2 KHz 
			end
			4'h1 :
			begin
				phase_inc = 32'h0003EEA2;//3 KHz
			end  
			4'h2 :
			begin
				phase_inc = 32'h00053E2D;//4 KHz
			end  
			4'h3 :
			begin
				phase_inc = 32'h00068DB8;//5 KHz
			end 
			4'h4 :
			begin
				phase_inc = 32'h0007DD44;//6 KHz
			end
			4'h5 :
			begin
				phase_inc = 32'h00092CCF;//7 KHz
			end  
			4'h6 :
			begin
				phase_inc = 32'h000A7C5A;//8 KHz
			end  
			4'h7 :
			begin
				phase_inc = 32'h000BCBE6;//9 KHz
			end
			4'h8 :
			begin
				phase_inc = 32'h000D1B71; //10 KHz center
			end
			4'h9 :
			begin
				phase_inc = 32'h000E6AFC;//11 KHz
			end  
			4'ha :
			begin
				phase_inc = 32'h000FBA88;//12 KHz
			end  
			4'hb :
			begin
				phase_inc = 32'h00110A13;//13 KHz
			end
			4'hc :
			begin
				phase_inc = 32'h0012599E;//14 KHz
			end
			4'hd :
			begin
				phase_inc = 32'h0013A92A;//15 KHz
			end  
			4'he :
			begin
				phase_inc = 32'h0014F8B5;//16 KHz
			end  
			4'hf :
			begin
				phase_inc = 32'h00164840;//17 KHz
			end    
		endcase

	end

endmodule

module freq_div (clk, clk_out);
	input clk;
	output clk_out;
	reg [1:0] r_reg =2'd 0;
	wire [1:0] r_nxt;
	reg clk_track = 0; 
	always @(posedge clk) 
	begin
		if (r_nxt == 2'b10)
		begin
			r_reg <= 2'd0;
			clk_track <= ~clk_track;
		end
		else 
			r_reg <= r_nxt;
		end
	assign r_nxt = r_reg + 2'd1;   	      
	assign clk_out = clk_track;
endmodule

module sincos_lut (
    input wire clk,
    input wire en,
    input wire [11:0] addr,
    output reg [11:0] sin_out,
    output reg [11:0] cos_out
);

// Define the size of the ROM
parameter ROM_SIZE = 4096;

// Define the ROMs as read-only memories
reg [11:0] SIN_ROM [0:ROM_SIZE-1];
reg [11:0] COS_ROM [0:ROM_SIZE-1];

// Initialize the ROM contents (replace with actual values)
//

// ROM select logic
always @(posedge clk) begin
    if (en) begin
        sin_out <= SIN_ROM[addr];
        cos_out <= COS_ROM[addr];
    end
end
//sin wave generated in matlab; converted from floating point to hex; and generated assignment code in python
	always@(posedge clk) begin

SIN_ROM[0] <= 12'h000; 
SIN_ROM[1] <= 12'h003; 
SIN_ROM[2] <= 12'h006; 
SIN_ROM[3] <= 12'h009; 
SIN_ROM[4] <= 12'h00d; 
SIN_ROM[5] <= 12'h010; 
SIN_ROM[6] <= 12'h013; 
SIN_ROM[7] <= 12'h016; 
SIN_ROM[8] <= 12'h019; 
SIN_ROM[9] <= 12'h01c; 
SIN_ROM[10] <= 12'h01f; 
SIN_ROM[11] <= 12'h023; 
SIN_ROM[12] <= 12'h026; 
SIN_ROM[13] <= 12'h029; 
SIN_ROM[14] <= 12'h02c; 
SIN_ROM[15] <= 12'h02f; 
SIN_ROM[16] <= 12'h032; 
SIN_ROM[17] <= 12'h035; 
SIN_ROM[18] <= 12'h039; 
SIN_ROM[19] <= 12'h03c; 
SIN_ROM[20] <= 12'h03f; 
SIN_ROM[21] <= 12'h042; 
SIN_ROM[22] <= 12'h045; 
SIN_ROM[23] <= 12'h048; 
SIN_ROM[24] <= 12'h04b; 
SIN_ROM[25] <= 12'h04e; 
SIN_ROM[26] <= 12'h052; 
SIN_ROM[27] <= 12'h055; 
SIN_ROM[28] <= 12'h058; 
SIN_ROM[29] <= 12'h05b; 
SIN_ROM[30] <= 12'h05e; 
SIN_ROM[31] <= 12'h061; 
SIN_ROM[32] <= 12'h064; 
SIN_ROM[33] <= 12'h068; 
SIN_ROM[34] <= 12'h06b; 
SIN_ROM[35] <= 12'h06e; 
SIN_ROM[36] <= 12'h071; 
SIN_ROM[37] <= 12'h074; 
SIN_ROM[38] <= 12'h077; 
SIN_ROM[39] <= 12'h07a; 
SIN_ROM[40] <= 12'h07e; 
SIN_ROM[41] <= 12'h081; 
SIN_ROM[42] <= 12'h084; 
SIN_ROM[43] <= 12'h087; 
SIN_ROM[44] <= 12'h08a; 
SIN_ROM[45] <= 12'h08d; 
SIN_ROM[46] <= 12'h090; 
SIN_ROM[47] <= 12'h093; 
SIN_ROM[48] <= 12'h097; 
SIN_ROM[49] <= 12'h09a; 
SIN_ROM[50] <= 12'h09d; 
SIN_ROM[51] <= 12'h0a0; 
SIN_ROM[52] <= 12'h0a3; 
SIN_ROM[53] <= 12'h0a6; 
SIN_ROM[54] <= 12'h0a9; 
SIN_ROM[55] <= 12'h0ac; 
SIN_ROM[56] <= 12'h0b0; 
SIN_ROM[57] <= 12'h0b3; 
SIN_ROM[58] <= 12'h0b6; 
SIN_ROM[59] <= 12'h0b9; 
SIN_ROM[60] <= 12'h0bc; 
SIN_ROM[61] <= 12'h0bf; 
SIN_ROM[62] <= 12'h0c2; 
SIN_ROM[63] <= 12'h0c6; 
SIN_ROM[64] <= 12'h0c9; 
SIN_ROM[65] <= 12'h0cc; 
SIN_ROM[66] <= 12'h0cf; 
SIN_ROM[67] <= 12'h0d2; 
SIN_ROM[68] <= 12'h0d5; 
SIN_ROM[69] <= 12'h0d8; 
SIN_ROM[70] <= 12'h0db; 
SIN_ROM[71] <= 12'h0df; 
SIN_ROM[72] <= 12'h0e2; 
SIN_ROM[73] <= 12'h0e5; 
SIN_ROM[74] <= 12'h0e8; 
SIN_ROM[75] <= 12'h0eb; 
SIN_ROM[76] <= 12'h0ee; 
SIN_ROM[77] <= 12'h0f1; 
SIN_ROM[78] <= 12'h0f4; 
SIN_ROM[79] <= 12'h0f7; 
SIN_ROM[80] <= 12'h0fb; 
SIN_ROM[81] <= 12'h0fe; 
SIN_ROM[82] <= 12'h101; 
SIN_ROM[83] <= 12'h104; 
SIN_ROM[84] <= 12'h107; 
SIN_ROM[85] <= 12'h10a; 
SIN_ROM[86] <= 12'h10d; 
SIN_ROM[87] <= 12'h110; 
SIN_ROM[88] <= 12'h113; 
SIN_ROM[89] <= 12'h117; 
SIN_ROM[90] <= 12'h11a; 
SIN_ROM[91] <= 12'h11d; 
SIN_ROM[92] <= 12'h120; 
SIN_ROM[93] <= 12'h123; 
SIN_ROM[94] <= 12'h126; 
SIN_ROM[95] <= 12'h129; 
SIN_ROM[96] <= 12'h12c; 
SIN_ROM[97] <= 12'h12f; 
SIN_ROM[98] <= 12'h133; 
SIN_ROM[99] <= 12'h136; 
SIN_ROM[100] <= 12'h139; 
SIN_ROM[101] <= 12'h13c; 
SIN_ROM[102] <= 12'h13f; 
SIN_ROM[103] <= 12'h142; 
SIN_ROM[104] <= 12'h145; 
SIN_ROM[105] <= 12'h148; 
SIN_ROM[106] <= 12'h14b; 
SIN_ROM[107] <= 12'h14e; 
SIN_ROM[108] <= 12'h152; 
SIN_ROM[109] <= 12'h155; 
SIN_ROM[110] <= 12'h158; 
SIN_ROM[111] <= 12'h15b; 
SIN_ROM[112] <= 12'h15e; 
SIN_ROM[113] <= 12'h161; 
SIN_ROM[114] <= 12'h164; 
SIN_ROM[115] <= 12'h167; 
SIN_ROM[116] <= 12'h16a; 
SIN_ROM[117] <= 12'h16d; 
SIN_ROM[118] <= 12'h171; 
SIN_ROM[119] <= 12'h174; 
SIN_ROM[120] <= 12'h177; 
SIN_ROM[121] <= 12'h17a; 
SIN_ROM[122] <= 12'h17d; 
SIN_ROM[123] <= 12'h180; 
SIN_ROM[124] <= 12'h183; 
SIN_ROM[125] <= 12'h186; 
SIN_ROM[126] <= 12'h189; 
SIN_ROM[127] <= 12'h18c; 
SIN_ROM[128] <= 12'h18f; 
SIN_ROM[129] <= 12'h192; 
SIN_ROM[130] <= 12'h196; 
SIN_ROM[131] <= 12'h199; 
SIN_ROM[132] <= 12'h19c; 
SIN_ROM[133] <= 12'h19f; 
SIN_ROM[134] <= 12'h1a2; 
SIN_ROM[135] <= 12'h1a5; 
SIN_ROM[136] <= 12'h1a8; 
SIN_ROM[137] <= 12'h1ab; 
SIN_ROM[138] <= 12'h1ae; 
SIN_ROM[139] <= 12'h1b1; 
SIN_ROM[140] <= 12'h1b4; 
SIN_ROM[141] <= 12'h1b7; 
SIN_ROM[142] <= 12'h1ba; 
SIN_ROM[143] <= 12'h1bd; 
SIN_ROM[144] <= 12'h1c1; 
SIN_ROM[145] <= 12'h1c4; 
SIN_ROM[146] <= 12'h1c7; 
SIN_ROM[147] <= 12'h1ca; 
SIN_ROM[148] <= 12'h1cd; 
SIN_ROM[149] <= 12'h1d0; 
SIN_ROM[150] <= 12'h1d3; 
SIN_ROM[151] <= 12'h1d6; 
SIN_ROM[152] <= 12'h1d9; 
SIN_ROM[153] <= 12'h1dc; 
SIN_ROM[154] <= 12'h1df; 
SIN_ROM[155] <= 12'h1e2; 
SIN_ROM[156] <= 12'h1e5; 
SIN_ROM[157] <= 12'h1e8; 
SIN_ROM[158] <= 12'h1eb; 
SIN_ROM[159] <= 12'h1ee; 
SIN_ROM[160] <= 12'h1f1; 
SIN_ROM[161] <= 12'h1f4; 
SIN_ROM[162] <= 12'h1f7; 
SIN_ROM[163] <= 12'h1fb; 
SIN_ROM[164] <= 12'h1fe; 
SIN_ROM[165] <= 12'h201; 
SIN_ROM[166] <= 12'h204; 
SIN_ROM[167] <= 12'h207; 
SIN_ROM[168] <= 12'h20a; 
SIN_ROM[169] <= 12'h20d; 
SIN_ROM[170] <= 12'h210; 
SIN_ROM[171] <= 12'h213; 
SIN_ROM[172] <= 12'h216; 
SIN_ROM[173] <= 12'h219; 
SIN_ROM[174] <= 12'h21c; 
SIN_ROM[175] <= 12'h21f; 
SIN_ROM[176] <= 12'h222; 
SIN_ROM[177] <= 12'h225; 
SIN_ROM[178] <= 12'h228; 
SIN_ROM[179] <= 12'h22b; 
SIN_ROM[180] <= 12'h22e; 
SIN_ROM[181] <= 12'h231; 
SIN_ROM[182] <= 12'h234; 
SIN_ROM[183] <= 12'h237; 
SIN_ROM[184] <= 12'h23a; 
SIN_ROM[185] <= 12'h23d; 
SIN_ROM[186] <= 12'h240; 
SIN_ROM[187] <= 12'h243; 
SIN_ROM[188] <= 12'h246; 
SIN_ROM[189] <= 12'h249; 
SIN_ROM[190] <= 12'h24c; 
SIN_ROM[191] <= 12'h24f; 
SIN_ROM[192] <= 12'h252; 
SIN_ROM[193] <= 12'h255; 
SIN_ROM[194] <= 12'h258; 
SIN_ROM[195] <= 12'h25b; 
SIN_ROM[196] <= 12'h25e; 
SIN_ROM[197] <= 12'h261; 
SIN_ROM[198] <= 12'h264; 
SIN_ROM[199] <= 12'h267; 
SIN_ROM[200] <= 12'h26a; 
SIN_ROM[201] <= 12'h26d; 
SIN_ROM[202] <= 12'h270; 
SIN_ROM[203] <= 12'h273; 
SIN_ROM[204] <= 12'h276; 
SIN_ROM[205] <= 12'h279; 
SIN_ROM[206] <= 12'h27c; 
SIN_ROM[207] <= 12'h27f; 
SIN_ROM[208] <= 12'h282; 
SIN_ROM[209] <= 12'h285; 
SIN_ROM[210] <= 12'h288; 
SIN_ROM[211] <= 12'h28b; 
SIN_ROM[212] <= 12'h28e; 
SIN_ROM[213] <= 12'h291; 
SIN_ROM[214] <= 12'h294; 
SIN_ROM[215] <= 12'h297; 
SIN_ROM[216] <= 12'h29a; 
SIN_ROM[217] <= 12'h29d; 
SIN_ROM[218] <= 12'h2a0; 
SIN_ROM[219] <= 12'h2a3; 
SIN_ROM[220] <= 12'h2a6; 
SIN_ROM[221] <= 12'h2a9; 
SIN_ROM[222] <= 12'h2ac; 
SIN_ROM[223] <= 12'h2af; 
SIN_ROM[224] <= 12'h2b2; 
SIN_ROM[225] <= 12'h2b5; 
SIN_ROM[226] <= 12'h2b8; 
SIN_ROM[227] <= 12'h2ba; 
SIN_ROM[228] <= 12'h2bd; 
SIN_ROM[229] <= 12'h2c0; 
SIN_ROM[230] <= 12'h2c3; 
SIN_ROM[231] <= 12'h2c6; 
SIN_ROM[232] <= 12'h2c9; 
SIN_ROM[233] <= 12'h2cc; 
SIN_ROM[234] <= 12'h2cf; 
SIN_ROM[235] <= 12'h2d2; 
SIN_ROM[236] <= 12'h2d5; 
SIN_ROM[237] <= 12'h2d8; 
SIN_ROM[238] <= 12'h2db; 
SIN_ROM[239] <= 12'h2de; 
SIN_ROM[240] <= 12'h2e1; 
SIN_ROM[241] <= 12'h2e4; 
SIN_ROM[242] <= 12'h2e7; 
SIN_ROM[243] <= 12'h2e9; 
SIN_ROM[244] <= 12'h2ec; 
SIN_ROM[245] <= 12'h2ef; 
SIN_ROM[246] <= 12'h2f2; 
SIN_ROM[247] <= 12'h2f5; 
SIN_ROM[248] <= 12'h2f8; 
SIN_ROM[249] <= 12'h2fb; 
SIN_ROM[250] <= 12'h2fe; 
SIN_ROM[251] <= 12'h301; 
SIN_ROM[252] <= 12'h304; 
SIN_ROM[253] <= 12'h307; 
SIN_ROM[254] <= 12'h30a; 
SIN_ROM[255] <= 12'h30c; 
SIN_ROM[256] <= 12'h30f; 
SIN_ROM[257] <= 12'h312; 
SIN_ROM[258] <= 12'h315; 
SIN_ROM[259] <= 12'h318; 
SIN_ROM[260] <= 12'h31b; 
SIN_ROM[261] <= 12'h31e; 
SIN_ROM[262] <= 12'h321; 
SIN_ROM[263] <= 12'h324; 
SIN_ROM[264] <= 12'h327; 
SIN_ROM[265] <= 12'h329; 
SIN_ROM[266] <= 12'h32c; 
SIN_ROM[267] <= 12'h32f; 
SIN_ROM[268] <= 12'h332; 
SIN_ROM[269] <= 12'h335; 
SIN_ROM[270] <= 12'h338; 
SIN_ROM[271] <= 12'h33b; 
SIN_ROM[272] <= 12'h33e; 
SIN_ROM[273] <= 12'h340; 
SIN_ROM[274] <= 12'h343; 
SIN_ROM[275] <= 12'h346; 
SIN_ROM[276] <= 12'h349; 
SIN_ROM[277] <= 12'h34c; 
SIN_ROM[278] <= 12'h34f; 
SIN_ROM[279] <= 12'h352; 
SIN_ROM[280] <= 12'h354; 
SIN_ROM[281] <= 12'h357; 
SIN_ROM[282] <= 12'h35a; 
SIN_ROM[283] <= 12'h35d; 
SIN_ROM[284] <= 12'h360; 
SIN_ROM[285] <= 12'h363; 
SIN_ROM[286] <= 12'h366; 
SIN_ROM[287] <= 12'h368; 
SIN_ROM[288] <= 12'h36b; 
SIN_ROM[289] <= 12'h36e; 
SIN_ROM[290] <= 12'h371; 
SIN_ROM[291] <= 12'h374; 
SIN_ROM[292] <= 12'h377; 
SIN_ROM[293] <= 12'h379; 
SIN_ROM[294] <= 12'h37c; 
SIN_ROM[295] <= 12'h37f; 
SIN_ROM[296] <= 12'h382; 
SIN_ROM[297] <= 12'h385; 
SIN_ROM[298] <= 12'h387; 
SIN_ROM[299] <= 12'h38a; 
SIN_ROM[300] <= 12'h38d; 
SIN_ROM[301] <= 12'h390; 
SIN_ROM[302] <= 12'h393; 
SIN_ROM[303] <= 12'h396; 
SIN_ROM[304] <= 12'h398; 
SIN_ROM[305] <= 12'h39b; 
SIN_ROM[306] <= 12'h39e; 
SIN_ROM[307] <= 12'h3a1; 
SIN_ROM[308] <= 12'h3a4; 
SIN_ROM[309] <= 12'h3a6; 
SIN_ROM[310] <= 12'h3a9; 
SIN_ROM[311] <= 12'h3ac; 
SIN_ROM[312] <= 12'h3af; 
SIN_ROM[313] <= 12'h3b2; 
SIN_ROM[314] <= 12'h3b4; 
SIN_ROM[315] <= 12'h3b7; 
SIN_ROM[316] <= 12'h3ba; 
SIN_ROM[317] <= 12'h3bd; 
SIN_ROM[318] <= 12'h3bf; 
SIN_ROM[319] <= 12'h3c2; 
SIN_ROM[320] <= 12'h3c5; 
SIN_ROM[321] <= 12'h3c8; 
SIN_ROM[322] <= 12'h3ca; 
SIN_ROM[323] <= 12'h3cd; 
SIN_ROM[324] <= 12'h3d0; 
SIN_ROM[325] <= 12'h3d3; 
SIN_ROM[326] <= 12'h3d6; 
SIN_ROM[327] <= 12'h3d8; 
SIN_ROM[328] <= 12'h3db; 
SIN_ROM[329] <= 12'h3de; 
SIN_ROM[330] <= 12'h3e1; 
SIN_ROM[331] <= 12'h3e3; 
SIN_ROM[332] <= 12'h3e6; 
SIN_ROM[333] <= 12'h3e9; 
SIN_ROM[334] <= 12'h3eb; 
SIN_ROM[335] <= 12'h3ee; 
SIN_ROM[336] <= 12'h3f1; 
SIN_ROM[337] <= 12'h3f4; 
SIN_ROM[338] <= 12'h3f6; 
SIN_ROM[339] <= 12'h3f9; 
SIN_ROM[340] <= 12'h3fc; 
SIN_ROM[341] <= 12'h3ff; 
SIN_ROM[342] <= 12'h401; 
SIN_ROM[343] <= 12'h404; 
SIN_ROM[344] <= 12'h407; 
SIN_ROM[345] <= 12'h409; 
SIN_ROM[346] <= 12'h40c; 
SIN_ROM[347] <= 12'h40f; 
SIN_ROM[348] <= 12'h412; 
SIN_ROM[349] <= 12'h414; 
SIN_ROM[350] <= 12'h417; 
SIN_ROM[351] <= 12'h41a; 
SIN_ROM[352] <= 12'h41c; 
SIN_ROM[353] <= 12'h41f; 
SIN_ROM[354] <= 12'h422; 
SIN_ROM[355] <= 12'h424; 
SIN_ROM[356] <= 12'h427; 
SIN_ROM[357] <= 12'h42a; 
SIN_ROM[358] <= 12'h42c; 
SIN_ROM[359] <= 12'h42f; 
SIN_ROM[360] <= 12'h432; 
SIN_ROM[361] <= 12'h435; 
SIN_ROM[362] <= 12'h437; 
SIN_ROM[363] <= 12'h43a; 
SIN_ROM[364] <= 12'h43d; 
SIN_ROM[365] <= 12'h43f; 
SIN_ROM[366] <= 12'h442; 
SIN_ROM[367] <= 12'h444; 
SIN_ROM[368] <= 12'h447; 
SIN_ROM[369] <= 12'h44a; 
SIN_ROM[370] <= 12'h44c; 
SIN_ROM[371] <= 12'h44f; 
SIN_ROM[372] <= 12'h452; 
SIN_ROM[373] <= 12'h454; 
SIN_ROM[374] <= 12'h457; 
SIN_ROM[375] <= 12'h45a; 
SIN_ROM[376] <= 12'h45c; 
SIN_ROM[377] <= 12'h45f; 
SIN_ROM[378] <= 12'h462; 
SIN_ROM[379] <= 12'h464; 
SIN_ROM[380] <= 12'h467; 
SIN_ROM[381] <= 12'h469; 
SIN_ROM[382] <= 12'h46c; 
SIN_ROM[383] <= 12'h46f; 
SIN_ROM[384] <= 12'h471; 
SIN_ROM[385] <= 12'h474; 
SIN_ROM[386] <= 12'h476; 
SIN_ROM[387] <= 12'h479; 
SIN_ROM[388] <= 12'h47c; 
SIN_ROM[389] <= 12'h47e; 
SIN_ROM[390] <= 12'h481; 
SIN_ROM[391] <= 12'h483; 
SIN_ROM[392] <= 12'h486; 
SIN_ROM[393] <= 12'h489; 
SIN_ROM[394] <= 12'h48b; 
SIN_ROM[395] <= 12'h48e; 
SIN_ROM[396] <= 12'h490; 
SIN_ROM[397] <= 12'h493; 
SIN_ROM[398] <= 12'h496; 
SIN_ROM[399] <= 12'h498; 
SIN_ROM[400] <= 12'h49b; 
SIN_ROM[401] <= 12'h49d; 
SIN_ROM[402] <= 12'h4a0; 
SIN_ROM[403] <= 12'h4a2; 
SIN_ROM[404] <= 12'h4a5; 
SIN_ROM[405] <= 12'h4a7; 
SIN_ROM[406] <= 12'h4aa; 
SIN_ROM[407] <= 12'h4ad; 
SIN_ROM[408] <= 12'h4af; 
SIN_ROM[409] <= 12'h4b2; 
SIN_ROM[410] <= 12'h4b4; 
SIN_ROM[411] <= 12'h4b7; 
SIN_ROM[412] <= 12'h4b9; 
SIN_ROM[413] <= 12'h4bc; 
SIN_ROM[414] <= 12'h4be; 
SIN_ROM[415] <= 12'h4c1; 
SIN_ROM[416] <= 12'h4c3; 
SIN_ROM[417] <= 12'h4c6; 
SIN_ROM[418] <= 12'h4c8; 
SIN_ROM[419] <= 12'h4cb; 
SIN_ROM[420] <= 12'h4cd; 
SIN_ROM[421] <= 12'h4d0; 
SIN_ROM[422] <= 12'h4d2; 
SIN_ROM[423] <= 12'h4d5; 
SIN_ROM[424] <= 12'h4d7; 
SIN_ROM[425] <= 12'h4da; 
SIN_ROM[426] <= 12'h4dc; 
SIN_ROM[427] <= 12'h4df; 
SIN_ROM[428] <= 12'h4e1; 
SIN_ROM[429] <= 12'h4e4; 
SIN_ROM[430] <= 12'h4e6; 
SIN_ROM[431] <= 12'h4e9; 
SIN_ROM[432] <= 12'h4eb; 
SIN_ROM[433] <= 12'h4ee; 
SIN_ROM[434] <= 12'h4f0; 
SIN_ROM[435] <= 12'h4f3; 
SIN_ROM[436] <= 12'h4f5; 
SIN_ROM[437] <= 12'h4f8; 
SIN_ROM[438] <= 12'h4fa; 
SIN_ROM[439] <= 12'h4fd; 
SIN_ROM[440] <= 12'h4ff; 
SIN_ROM[441] <= 12'h502; 
SIN_ROM[442] <= 12'h504; 
SIN_ROM[443] <= 12'h506; 
SIN_ROM[444] <= 12'h509; 
SIN_ROM[445] <= 12'h50b; 
SIN_ROM[446] <= 12'h50e; 
SIN_ROM[447] <= 12'h510; 
SIN_ROM[448] <= 12'h513; 
SIN_ROM[449] <= 12'h515; 
SIN_ROM[450] <= 12'h517; 
SIN_ROM[451] <= 12'h51a; 
SIN_ROM[452] <= 12'h51c; 
SIN_ROM[453] <= 12'h51f; 
SIN_ROM[454] <= 12'h521; 
SIN_ROM[455] <= 12'h524; 
SIN_ROM[456] <= 12'h526; 
SIN_ROM[457] <= 12'h528; 
SIN_ROM[458] <= 12'h52b; 
SIN_ROM[459] <= 12'h52d; 
SIN_ROM[460] <= 12'h530; 
SIN_ROM[461] <= 12'h532; 
SIN_ROM[462] <= 12'h534; 
SIN_ROM[463] <= 12'h537; 
SIN_ROM[464] <= 12'h539; 
SIN_ROM[465] <= 12'h53b; 
SIN_ROM[466] <= 12'h53e; 
SIN_ROM[467] <= 12'h540; 
SIN_ROM[468] <= 12'h543; 
SIN_ROM[469] <= 12'h545; 
SIN_ROM[470] <= 12'h547; 
SIN_ROM[471] <= 12'h54a; 
SIN_ROM[472] <= 12'h54c; 
SIN_ROM[473] <= 12'h54e; 
SIN_ROM[474] <= 12'h551; 
SIN_ROM[475] <= 12'h553; 
SIN_ROM[476] <= 12'h555; 
SIN_ROM[477] <= 12'h558; 
SIN_ROM[478] <= 12'h55a; 
SIN_ROM[479] <= 12'h55c; 
SIN_ROM[480] <= 12'h55f; 
SIN_ROM[481] <= 12'h561; 
SIN_ROM[482] <= 12'h563; 
SIN_ROM[483] <= 12'h566; 
SIN_ROM[484] <= 12'h568; 
SIN_ROM[485] <= 12'h56a; 
SIN_ROM[486] <= 12'h56d; 
SIN_ROM[487] <= 12'h56f; 
SIN_ROM[488] <= 12'h571; 
SIN_ROM[489] <= 12'h573; 
SIN_ROM[490] <= 12'h576; 
SIN_ROM[491] <= 12'h578; 
SIN_ROM[492] <= 12'h57a; 
SIN_ROM[493] <= 12'h57d; 
SIN_ROM[494] <= 12'h57f; 
SIN_ROM[495] <= 12'h581; 
SIN_ROM[496] <= 12'h583; 
SIN_ROM[497] <= 12'h586; 
SIN_ROM[498] <= 12'h588; 
SIN_ROM[499] <= 12'h58a; 
SIN_ROM[500] <= 12'h58d; 
SIN_ROM[501] <= 12'h58f; 
SIN_ROM[502] <= 12'h591; 
SIN_ROM[503] <= 12'h593; 
SIN_ROM[504] <= 12'h596; 
SIN_ROM[505] <= 12'h598; 
SIN_ROM[506] <= 12'h59a; 
SIN_ROM[507] <= 12'h59c; 
SIN_ROM[508] <= 12'h59f; 
SIN_ROM[509] <= 12'h5a1; 
SIN_ROM[510] <= 12'h5a3; 
SIN_ROM[511] <= 12'h5a5; 
SIN_ROM[512] <= 12'h5a7; 
SIN_ROM[513] <= 12'h5aa; 
SIN_ROM[514] <= 12'h5ac; 
SIN_ROM[515] <= 12'h5ae; 
SIN_ROM[516] <= 12'h5b0; 
SIN_ROM[517] <= 12'h5b3; 
SIN_ROM[518] <= 12'h5b5; 
SIN_ROM[519] <= 12'h5b7; 
SIN_ROM[520] <= 12'h5b9; 
SIN_ROM[521] <= 12'h5bb; 
SIN_ROM[522] <= 12'h5bd; 
SIN_ROM[523] <= 12'h5c0; 
SIN_ROM[524] <= 12'h5c2; 
SIN_ROM[525] <= 12'h5c4; 
SIN_ROM[526] <= 12'h5c6; 
SIN_ROM[527] <= 12'h5c8; 
SIN_ROM[528] <= 12'h5cb; 
SIN_ROM[529] <= 12'h5cd; 
SIN_ROM[530] <= 12'h5cf; 
SIN_ROM[531] <= 12'h5d1; 
SIN_ROM[532] <= 12'h5d3; 
SIN_ROM[533] <= 12'h5d5; 
SIN_ROM[534] <= 12'h5d7; 
SIN_ROM[535] <= 12'h5da; 
SIN_ROM[536] <= 12'h5dc; 
SIN_ROM[537] <= 12'h5de; 
SIN_ROM[538] <= 12'h5e0; 
SIN_ROM[539] <= 12'h5e2; 
SIN_ROM[540] <= 12'h5e4; 
SIN_ROM[541] <= 12'h5e6; 
SIN_ROM[542] <= 12'h5e9; 
SIN_ROM[543] <= 12'h5eb; 
SIN_ROM[544] <= 12'h5ed; 
SIN_ROM[545] <= 12'h5ef; 
SIN_ROM[546] <= 12'h5f1; 
SIN_ROM[547] <= 12'h5f3; 
SIN_ROM[548] <= 12'h5f5; 
SIN_ROM[549] <= 12'h5f7; 
SIN_ROM[550] <= 12'h5f9; 
SIN_ROM[551] <= 12'h5fb; 
SIN_ROM[552] <= 12'h5fd; 
SIN_ROM[553] <= 12'h600; 
SIN_ROM[554] <= 12'h602; 
SIN_ROM[555] <= 12'h604; 
SIN_ROM[556] <= 12'h606; 
SIN_ROM[557] <= 12'h608; 
SIN_ROM[558] <= 12'h60a; 
SIN_ROM[559] <= 12'h60c; 
SIN_ROM[560] <= 12'h60e; 
SIN_ROM[561] <= 12'h610; 
SIN_ROM[562] <= 12'h612; 
SIN_ROM[563] <= 12'h614; 
SIN_ROM[564] <= 12'h616; 
SIN_ROM[565] <= 12'h618; 
SIN_ROM[566] <= 12'h61a; 
SIN_ROM[567] <= 12'h61c; 
SIN_ROM[568] <= 12'h61e; 
SIN_ROM[569] <= 12'h620; 
SIN_ROM[570] <= 12'h622; 
SIN_ROM[571] <= 12'h624; 
SIN_ROM[572] <= 12'h626; 
SIN_ROM[573] <= 12'h628; 
SIN_ROM[574] <= 12'h62a; 
SIN_ROM[575] <= 12'h62c; 
SIN_ROM[576] <= 12'h62e; 
SIN_ROM[577] <= 12'h630; 
SIN_ROM[578] <= 12'h632; 
SIN_ROM[579] <= 12'h634; 
SIN_ROM[580] <= 12'h636; 
SIN_ROM[581] <= 12'h638; 
SIN_ROM[582] <= 12'h63a; 
SIN_ROM[583] <= 12'h63c; 
SIN_ROM[584] <= 12'h63e; 
SIN_ROM[585] <= 12'h640; 
SIN_ROM[586] <= 12'h642; 
SIN_ROM[587] <= 12'h644; 
SIN_ROM[588] <= 12'h646; 
SIN_ROM[589] <= 12'h648; 
SIN_ROM[590] <= 12'h64a; 
SIN_ROM[591] <= 12'h64c; 
SIN_ROM[592] <= 12'h64e; 
SIN_ROM[593] <= 12'h650; 
SIN_ROM[594] <= 12'h652; 
SIN_ROM[595] <= 12'h654; 
SIN_ROM[596] <= 12'h655; 
SIN_ROM[597] <= 12'h657; 
SIN_ROM[598] <= 12'h659; 
SIN_ROM[599] <= 12'h65b; 
SIN_ROM[600] <= 12'h65d; 
SIN_ROM[601] <= 12'h65f; 
SIN_ROM[602] <= 12'h661; 
SIN_ROM[603] <= 12'h663; 
SIN_ROM[604] <= 12'h665; 
SIN_ROM[605] <= 12'h667; 
SIN_ROM[606] <= 12'h668; 
SIN_ROM[607] <= 12'h66a; 
SIN_ROM[608] <= 12'h66c; 
SIN_ROM[609] <= 12'h66e; 
SIN_ROM[610] <= 12'h670; 
SIN_ROM[611] <= 12'h672; 
SIN_ROM[612] <= 12'h674; 
SIN_ROM[613] <= 12'h675; 
SIN_ROM[614] <= 12'h677; 
SIN_ROM[615] <= 12'h679; 
SIN_ROM[616] <= 12'h67b; 
SIN_ROM[617] <= 12'h67d; 
SIN_ROM[618] <= 12'h67f; 
SIN_ROM[619] <= 12'h681; 
SIN_ROM[620] <= 12'h682; 
SIN_ROM[621] <= 12'h684; 
SIN_ROM[622] <= 12'h686; 
SIN_ROM[623] <= 12'h688; 
SIN_ROM[624] <= 12'h68a; 
SIN_ROM[625] <= 12'h68b; 
SIN_ROM[626] <= 12'h68d; 
SIN_ROM[627] <= 12'h68f; 
SIN_ROM[628] <= 12'h691; 
SIN_ROM[629] <= 12'h693; 
SIN_ROM[630] <= 12'h694; 
SIN_ROM[631] <= 12'h696; 
SIN_ROM[632] <= 12'h698; 
SIN_ROM[633] <= 12'h69a; 
SIN_ROM[634] <= 12'h69b; 
SIN_ROM[635] <= 12'h69d; 
SIN_ROM[636] <= 12'h69f; 
SIN_ROM[637] <= 12'h6a1; 
SIN_ROM[638] <= 12'h6a3; 
SIN_ROM[639] <= 12'h6a4; 
SIN_ROM[640] <= 12'h6a6; 
SIN_ROM[641] <= 12'h6a8; 
SIN_ROM[642] <= 12'h6a9; 
SIN_ROM[643] <= 12'h6ab; 
SIN_ROM[644] <= 12'h6ad; 
SIN_ROM[645] <= 12'h6af; 
SIN_ROM[646] <= 12'h6b0; 
SIN_ROM[647] <= 12'h6b2; 
SIN_ROM[648] <= 12'h6b4; 
SIN_ROM[649] <= 12'h6b6; 
SIN_ROM[650] <= 12'h6b7; 
SIN_ROM[651] <= 12'h6b9; 
SIN_ROM[652] <= 12'h6bb; 
SIN_ROM[653] <= 12'h6bc; 
SIN_ROM[654] <= 12'h6be; 
SIN_ROM[655] <= 12'h6c0; 
SIN_ROM[656] <= 12'h6c1; 
SIN_ROM[657] <= 12'h6c3; 
SIN_ROM[658] <= 12'h6c5; 
SIN_ROM[659] <= 12'h6c6; 
SIN_ROM[660] <= 12'h6c8; 
SIN_ROM[661] <= 12'h6ca; 
SIN_ROM[662] <= 12'h6cb; 
SIN_ROM[663] <= 12'h6cd; 
SIN_ROM[664] <= 12'h6cf; 
SIN_ROM[665] <= 12'h6d0; 
SIN_ROM[666] <= 12'h6d2; 
SIN_ROM[667] <= 12'h6d4; 
SIN_ROM[668] <= 12'h6d5; 
SIN_ROM[669] <= 12'h6d7; 
SIN_ROM[670] <= 12'h6d9; 
SIN_ROM[671] <= 12'h6da; 
SIN_ROM[672] <= 12'h6dc; 
SIN_ROM[673] <= 12'h6dd; 
SIN_ROM[674] <= 12'h6df; 
SIN_ROM[675] <= 12'h6e1; 
SIN_ROM[676] <= 12'h6e2; 
SIN_ROM[677] <= 12'h6e4; 
SIN_ROM[678] <= 12'h6e5; 
SIN_ROM[679] <= 12'h6e7; 
SIN_ROM[680] <= 12'h6e9; 
SIN_ROM[681] <= 12'h6ea; 
SIN_ROM[682] <= 12'h6ec; 
SIN_ROM[683] <= 12'h6ed; 
SIN_ROM[684] <= 12'h6ef; 
SIN_ROM[685] <= 12'h6f0; 
SIN_ROM[686] <= 12'h6f2; 
SIN_ROM[687] <= 12'h6f4; 
SIN_ROM[688] <= 12'h6f5; 
SIN_ROM[689] <= 12'h6f7; 
SIN_ROM[690] <= 12'h6f8; 
SIN_ROM[691] <= 12'h6fa; 
SIN_ROM[692] <= 12'h6fb; 
SIN_ROM[693] <= 12'h6fd; 
SIN_ROM[694] <= 12'h6fe; 
SIN_ROM[695] <= 12'h700; 
SIN_ROM[696] <= 12'h701; 
SIN_ROM[697] <= 12'h703; 
SIN_ROM[698] <= 12'h704; 
SIN_ROM[699] <= 12'h706; 
SIN_ROM[700] <= 12'h707; 
SIN_ROM[701] <= 12'h709; 
SIN_ROM[702] <= 12'h70a; 
SIN_ROM[703] <= 12'h70c; 
SIN_ROM[704] <= 12'h70d; 
SIN_ROM[705] <= 12'h70f; 
SIN_ROM[706] <= 12'h710; 
SIN_ROM[707] <= 12'h712; 
SIN_ROM[708] <= 12'h713; 
SIN_ROM[709] <= 12'h715; 
SIN_ROM[710] <= 12'h716; 
SIN_ROM[711] <= 12'h718; 
SIN_ROM[712] <= 12'h719; 
SIN_ROM[713] <= 12'h71a; 
SIN_ROM[714] <= 12'h71c; 
SIN_ROM[715] <= 12'h71d; 
SIN_ROM[716] <= 12'h71f; 
SIN_ROM[717] <= 12'h720; 
SIN_ROM[718] <= 12'h722; 
SIN_ROM[719] <= 12'h723; 
SIN_ROM[720] <= 12'h724; 
SIN_ROM[721] <= 12'h726; 
SIN_ROM[722] <= 12'h727; 
SIN_ROM[723] <= 12'h729; 
SIN_ROM[724] <= 12'h72a; 
SIN_ROM[725] <= 12'h72b; 
SIN_ROM[726] <= 12'h72d; 
SIN_ROM[727] <= 12'h72e; 
SIN_ROM[728] <= 12'h730; 
SIN_ROM[729] <= 12'h731; 
SIN_ROM[730] <= 12'h732; 
SIN_ROM[731] <= 12'h734; 
SIN_ROM[732] <= 12'h735; 
SIN_ROM[733] <= 12'h736; 
SIN_ROM[734] <= 12'h738; 
SIN_ROM[735] <= 12'h739; 
SIN_ROM[736] <= 12'h73a; 
SIN_ROM[737] <= 12'h73c; 
SIN_ROM[738] <= 12'h73d; 
SIN_ROM[739] <= 12'h73e; 
SIN_ROM[740] <= 12'h740; 
SIN_ROM[741] <= 12'h741; 
SIN_ROM[742] <= 12'h742; 
SIN_ROM[743] <= 12'h744; 
SIN_ROM[744] <= 12'h745; 
SIN_ROM[745] <= 12'h746; 
SIN_ROM[746] <= 12'h748; 
SIN_ROM[747] <= 12'h749; 
SIN_ROM[748] <= 12'h74a; 
SIN_ROM[749] <= 12'h74c; 
SIN_ROM[750] <= 12'h74d; 
SIN_ROM[751] <= 12'h74e; 
SIN_ROM[752] <= 12'h74f; 
SIN_ROM[753] <= 12'h751; 
SIN_ROM[754] <= 12'h752; 
SIN_ROM[755] <= 12'h753; 
SIN_ROM[756] <= 12'h754; 
SIN_ROM[757] <= 12'h756; 
SIN_ROM[758] <= 12'h757; 
SIN_ROM[759] <= 12'h758; 
SIN_ROM[760] <= 12'h759; 
SIN_ROM[761] <= 12'h75b; 
SIN_ROM[762] <= 12'h75c; 
SIN_ROM[763] <= 12'h75d; 
SIN_ROM[764] <= 12'h75e; 
SIN_ROM[765] <= 12'h760; 
SIN_ROM[766] <= 12'h761; 
SIN_ROM[767] <= 12'h762; 
SIN_ROM[768] <= 12'h763; 
SIN_ROM[769] <= 12'h764; 
SIN_ROM[770] <= 12'h766; 
SIN_ROM[771] <= 12'h767; 
SIN_ROM[772] <= 12'h768; 
SIN_ROM[773] <= 12'h769; 
SIN_ROM[774] <= 12'h76a; 
SIN_ROM[775] <= 12'h76b; 
SIN_ROM[776] <= 12'h76d; 
SIN_ROM[777] <= 12'h76e; 
SIN_ROM[778] <= 12'h76f; 
SIN_ROM[779] <= 12'h770; 
SIN_ROM[780] <= 12'h771; 
SIN_ROM[781] <= 12'h772; 
SIN_ROM[782] <= 12'h774; 
SIN_ROM[783] <= 12'h775; 
SIN_ROM[784] <= 12'h776; 
SIN_ROM[785] <= 12'h777; 
SIN_ROM[786] <= 12'h778; 
SIN_ROM[787] <= 12'h779; 
SIN_ROM[788] <= 12'h77a; 
SIN_ROM[789] <= 12'h77b; 
SIN_ROM[790] <= 12'h77d; 
SIN_ROM[791] <= 12'h77e; 
SIN_ROM[792] <= 12'h77f; 
SIN_ROM[793] <= 12'h780; 
SIN_ROM[794] <= 12'h781; 
SIN_ROM[795] <= 12'h782; 
SIN_ROM[796] <= 12'h783; 
SIN_ROM[797] <= 12'h784; 
SIN_ROM[798] <= 12'h785; 
SIN_ROM[799] <= 12'h786; 
SIN_ROM[800] <= 12'h787; 
SIN_ROM[801] <= 12'h788; 
SIN_ROM[802] <= 12'h789; 
SIN_ROM[803] <= 12'h78a; 
SIN_ROM[804] <= 12'h78c; 
SIN_ROM[805] <= 12'h78d; 
SIN_ROM[806] <= 12'h78e; 
SIN_ROM[807] <= 12'h78f; 
SIN_ROM[808] <= 12'h790; 
SIN_ROM[809] <= 12'h791; 
SIN_ROM[810] <= 12'h792; 
SIN_ROM[811] <= 12'h793; 
SIN_ROM[812] <= 12'h794; 
SIN_ROM[813] <= 12'h795; 
SIN_ROM[814] <= 12'h796; 
SIN_ROM[815] <= 12'h797; 
SIN_ROM[816] <= 12'h798; 
SIN_ROM[817] <= 12'h799; 
SIN_ROM[818] <= 12'h79a; 
SIN_ROM[819] <= 12'h79b; 
SIN_ROM[820] <= 12'h79c; 
SIN_ROM[821] <= 12'h79d; 
SIN_ROM[822] <= 12'h79e; 
SIN_ROM[823] <= 12'h79e; 
SIN_ROM[824] <= 12'h79f; 
SIN_ROM[825] <= 12'h7a0; 
SIN_ROM[826] <= 12'h7a1; 
SIN_ROM[827] <= 12'h7a2; 
SIN_ROM[828] <= 12'h7a3; 
SIN_ROM[829] <= 12'h7a4; 
SIN_ROM[830] <= 12'h7a5; 
SIN_ROM[831] <= 12'h7a6; 
SIN_ROM[832] <= 12'h7a7; 
SIN_ROM[833] <= 12'h7a8; 
SIN_ROM[834] <= 12'h7a9; 
SIN_ROM[835] <= 12'h7aa; 
SIN_ROM[836] <= 12'h7aa; 
SIN_ROM[837] <= 12'h7ab; 
SIN_ROM[838] <= 12'h7ac; 
SIN_ROM[839] <= 12'h7ad; 
SIN_ROM[840] <= 12'h7ae; 
SIN_ROM[841] <= 12'h7af; 
SIN_ROM[842] <= 12'h7b0; 
SIN_ROM[843] <= 12'h7b1; 
SIN_ROM[844] <= 12'h7b1; 
SIN_ROM[845] <= 12'h7b2; 
SIN_ROM[846] <= 12'h7b3; 
SIN_ROM[847] <= 12'h7b4; 
SIN_ROM[848] <= 12'h7b5; 
SIN_ROM[849] <= 12'h7b6; 
SIN_ROM[850] <= 12'h7b7; 
SIN_ROM[851] <= 12'h7b7; 
SIN_ROM[852] <= 12'h7b8; 
SIN_ROM[853] <= 12'h7b9; 
SIN_ROM[854] <= 12'h7ba; 
SIN_ROM[855] <= 12'h7bb; 
SIN_ROM[856] <= 12'h7bb; 
SIN_ROM[857] <= 12'h7bc; 
SIN_ROM[858] <= 12'h7bd; 
SIN_ROM[859] <= 12'h7be; 
SIN_ROM[860] <= 12'h7bf; 
SIN_ROM[861] <= 12'h7bf; 
SIN_ROM[862] <= 12'h7c0; 
SIN_ROM[863] <= 12'h7c1; 
SIN_ROM[864] <= 12'h7c2; 
SIN_ROM[865] <= 12'h7c2; 
SIN_ROM[866] <= 12'h7c3; 
SIN_ROM[867] <= 12'h7c4; 
SIN_ROM[868] <= 12'h7c5; 
SIN_ROM[869] <= 12'h7c5; 
SIN_ROM[870] <= 12'h7c6; 
SIN_ROM[871] <= 12'h7c7; 
SIN_ROM[872] <= 12'h7c8; 
SIN_ROM[873] <= 12'h7c8; 
SIN_ROM[874] <= 12'h7c9; 
SIN_ROM[875] <= 12'h7ca; 
SIN_ROM[876] <= 12'h7ca; 
SIN_ROM[877] <= 12'h7cb; 
SIN_ROM[878] <= 12'h7cc; 
SIN_ROM[879] <= 12'h7cd; 
SIN_ROM[880] <= 12'h7cd; 
SIN_ROM[881] <= 12'h7ce; 
SIN_ROM[882] <= 12'h7cf; 
SIN_ROM[883] <= 12'h7cf; 
SIN_ROM[884] <= 12'h7d0; 
SIN_ROM[885] <= 12'h7d1; 
SIN_ROM[886] <= 12'h7d1; 
SIN_ROM[887] <= 12'h7d2; 
SIN_ROM[888] <= 12'h7d3; 
SIN_ROM[889] <= 12'h7d3; 
SIN_ROM[890] <= 12'h7d4; 
SIN_ROM[891] <= 12'h7d5; 
SIN_ROM[892] <= 12'h7d5; 
SIN_ROM[893] <= 12'h7d6; 
SIN_ROM[894] <= 12'h7d6; 
SIN_ROM[895] <= 12'h7d7; 
SIN_ROM[896] <= 12'h7d8; 
SIN_ROM[897] <= 12'h7d8; 
SIN_ROM[898] <= 12'h7d9; 
SIN_ROM[899] <= 12'h7d9; 
SIN_ROM[900] <= 12'h7da; 
SIN_ROM[901] <= 12'h7db; 
SIN_ROM[902] <= 12'h7db; 
SIN_ROM[903] <= 12'h7dc; 
SIN_ROM[904] <= 12'h7dc; 
SIN_ROM[905] <= 12'h7dd; 
SIN_ROM[906] <= 12'h7de; 
SIN_ROM[907] <= 12'h7de; 
SIN_ROM[908] <= 12'h7df; 
SIN_ROM[909] <= 12'h7df; 
SIN_ROM[910] <= 12'h7e0; 
SIN_ROM[911] <= 12'h7e0; 
SIN_ROM[912] <= 12'h7e1; 
SIN_ROM[913] <= 12'h7e1; 
SIN_ROM[914] <= 12'h7e2; 
SIN_ROM[915] <= 12'h7e2; 
SIN_ROM[916] <= 12'h7e3; 
SIN_ROM[917] <= 12'h7e3; 
SIN_ROM[918] <= 12'h7e4; 
SIN_ROM[919] <= 12'h7e5; 
SIN_ROM[920] <= 12'h7e5; 
SIN_ROM[921] <= 12'h7e6; 
SIN_ROM[922] <= 12'h7e6; 
SIN_ROM[923] <= 12'h7e6; 
SIN_ROM[924] <= 12'h7e7; 
SIN_ROM[925] <= 12'h7e7; 
SIN_ROM[926] <= 12'h7e8; 
SIN_ROM[927] <= 12'h7e8; 
SIN_ROM[928] <= 12'h7e9; 
SIN_ROM[929] <= 12'h7e9; 
SIN_ROM[930] <= 12'h7ea; 
SIN_ROM[931] <= 12'h7ea; 
SIN_ROM[932] <= 12'h7eb; 
SIN_ROM[933] <= 12'h7eb; 
SIN_ROM[934] <= 12'h7ec; 
SIN_ROM[935] <= 12'h7ec; 
SIN_ROM[936] <= 12'h7ec; 
SIN_ROM[937] <= 12'h7ed; 
SIN_ROM[938] <= 12'h7ed; 
SIN_ROM[939] <= 12'h7ee; 
SIN_ROM[940] <= 12'h7ee; 
SIN_ROM[941] <= 12'h7ee; 
SIN_ROM[942] <= 12'h7ef; 
SIN_ROM[943] <= 12'h7ef; 
SIN_ROM[944] <= 12'h7f0; 
SIN_ROM[945] <= 12'h7f0; 
SIN_ROM[946] <= 12'h7f0; 
SIN_ROM[947] <= 12'h7f1; 
SIN_ROM[948] <= 12'h7f1; 
SIN_ROM[949] <= 12'h7f1; 
SIN_ROM[950] <= 12'h7f2; 
SIN_ROM[951] <= 12'h7f2; 
SIN_ROM[952] <= 12'h7f3; 
SIN_ROM[953] <= 12'h7f3; 
SIN_ROM[954] <= 12'h7f3; 
SIN_ROM[955] <= 12'h7f4; 
SIN_ROM[956] <= 12'h7f4; 
SIN_ROM[957] <= 12'h7f4; 
SIN_ROM[958] <= 12'h7f5; 
SIN_ROM[959] <= 12'h7f5; 
SIN_ROM[960] <= 12'h7f5; 
SIN_ROM[961] <= 12'h7f5; 
SIN_ROM[962] <= 12'h7f6; 
SIN_ROM[963] <= 12'h7f6; 
SIN_ROM[964] <= 12'h7f6; 
SIN_ROM[965] <= 12'h7f7; 
SIN_ROM[966] <= 12'h7f7; 
SIN_ROM[967] <= 12'h7f7; 
SIN_ROM[968] <= 12'h7f7; 
SIN_ROM[969] <= 12'h7f8; 
SIN_ROM[970] <= 12'h7f8; 
SIN_ROM[971] <= 12'h7f8; 
SIN_ROM[972] <= 12'h7f8; 
SIN_ROM[973] <= 12'h7f9; 
SIN_ROM[974] <= 12'h7f9; 
SIN_ROM[975] <= 12'h7f9; 
SIN_ROM[976] <= 12'h7f9; 
SIN_ROM[977] <= 12'h7fa; 
SIN_ROM[978] <= 12'h7fa; 
SIN_ROM[979] <= 12'h7fa; 
SIN_ROM[980] <= 12'h7fa; 
SIN_ROM[981] <= 12'h7fb; 
SIN_ROM[982] <= 12'h7fb; 
SIN_ROM[983] <= 12'h7fb; 
SIN_ROM[984] <= 12'h7fb; 
SIN_ROM[985] <= 12'h7fb; 
SIN_ROM[986] <= 12'h7fc; 
SIN_ROM[987] <= 12'h7fc; 
SIN_ROM[988] <= 12'h7fc; 
SIN_ROM[989] <= 12'h7fc; 
SIN_ROM[990] <= 12'h7fc; 
SIN_ROM[991] <= 12'h7fc; 
SIN_ROM[992] <= 12'h7fd; 
SIN_ROM[993] <= 12'h7fd; 
SIN_ROM[994] <= 12'h7fd; 
SIN_ROM[995] <= 12'h7fd; 
SIN_ROM[996] <= 12'h7fd; 
SIN_ROM[997] <= 12'h7fd; 
SIN_ROM[998] <= 12'h7fd; 
SIN_ROM[999] <= 12'h7fd; 
SIN_ROM[1000] <= 12'h7fe; 
SIN_ROM[1001] <= 12'h7fe; 
SIN_ROM[1002] <= 12'h7fe; 
SIN_ROM[1003] <= 12'h7fe; 
SIN_ROM[1004] <= 12'h7fe; 
SIN_ROM[1005] <= 12'h7fe; 
SIN_ROM[1006] <= 12'h7fe; 
SIN_ROM[1007] <= 12'h7fe; 
SIN_ROM[1008] <= 12'h7fe; 
SIN_ROM[1009] <= 12'h7fe; 
SIN_ROM[1010] <= 12'h7ff; 
SIN_ROM[1011] <= 12'h7ff; 
SIN_ROM[1012] <= 12'h7ff; 
SIN_ROM[1013] <= 12'h7ff; 
SIN_ROM[1014] <= 12'h7ff; 
SIN_ROM[1015] <= 12'h7ff; 
SIN_ROM[1016] <= 12'h7ff; 
SIN_ROM[1017] <= 12'h7ff; 
SIN_ROM[1018] <= 12'h7ff; 
SIN_ROM[1019] <= 12'h7ff; 
SIN_ROM[1020] <= 12'h7ff; 
SIN_ROM[1021] <= 12'h7ff; 
SIN_ROM[1022] <= 12'h7ff; 
SIN_ROM[1023] <= 12'h7ff; 
SIN_ROM[1024] <= 12'h7ff; 
SIN_ROM[1025] <= 12'h7ff; 
SIN_ROM[1026] <= 12'h7ff; 
SIN_ROM[1027] <= 12'h7ff; 
SIN_ROM[1028] <= 12'h7ff; 
SIN_ROM[1029] <= 12'h7ff; 
SIN_ROM[1030] <= 12'h7ff; 
SIN_ROM[1031] <= 12'h7ff; 
SIN_ROM[1032] <= 12'h7ff; 
SIN_ROM[1033] <= 12'h7ff; 
SIN_ROM[1034] <= 12'h7ff; 
SIN_ROM[1035] <= 12'h7ff; 
SIN_ROM[1036] <= 12'h7ff; 
SIN_ROM[1037] <= 12'h7ff; 
SIN_ROM[1038] <= 12'h7ff; 
SIN_ROM[1039] <= 12'h7fe; 
SIN_ROM[1040] <= 12'h7fe; 
SIN_ROM[1041] <= 12'h7fe; 
SIN_ROM[1042] <= 12'h7fe; 
SIN_ROM[1043] <= 12'h7fe; 
SIN_ROM[1044] <= 12'h7fe; 
SIN_ROM[1045] <= 12'h7fe; 
SIN_ROM[1046] <= 12'h7fe; 
SIN_ROM[1047] <= 12'h7fe; 
SIN_ROM[1048] <= 12'h7fe; 
SIN_ROM[1049] <= 12'h7fd; 
SIN_ROM[1050] <= 12'h7fd; 
SIN_ROM[1051] <= 12'h7fd; 
SIN_ROM[1052] <= 12'h7fd; 
SIN_ROM[1053] <= 12'h7fd; 
SIN_ROM[1054] <= 12'h7fd; 
SIN_ROM[1055] <= 12'h7fd; 
SIN_ROM[1056] <= 12'h7fd; 
SIN_ROM[1057] <= 12'h7fc; 
SIN_ROM[1058] <= 12'h7fc; 
SIN_ROM[1059] <= 12'h7fc; 
SIN_ROM[1060] <= 12'h7fc; 
SIN_ROM[1061] <= 12'h7fc; 
SIN_ROM[1062] <= 12'h7fc; 
SIN_ROM[1063] <= 12'h7fb; 
SIN_ROM[1064] <= 12'h7fb; 
SIN_ROM[1065] <= 12'h7fb; 
SIN_ROM[1066] <= 12'h7fb; 
SIN_ROM[1067] <= 12'h7fb; 
SIN_ROM[1068] <= 12'h7fa; 
SIN_ROM[1069] <= 12'h7fa; 
SIN_ROM[1070] <= 12'h7fa; 
SIN_ROM[1071] <= 12'h7fa; 
SIN_ROM[1072] <= 12'h7f9; 
SIN_ROM[1073] <= 12'h7f9; 
SIN_ROM[1074] <= 12'h7f9; 
SIN_ROM[1075] <= 12'h7f9; 
SIN_ROM[1076] <= 12'h7f8; 
SIN_ROM[1077] <= 12'h7f8; 
SIN_ROM[1078] <= 12'h7f8; 
SIN_ROM[1079] <= 12'h7f8; 
SIN_ROM[1080] <= 12'h7f7; 
SIN_ROM[1081] <= 12'h7f7; 
SIN_ROM[1082] <= 12'h7f7; 
SIN_ROM[1083] <= 12'h7f7; 
SIN_ROM[1084] <= 12'h7f6; 
SIN_ROM[1085] <= 12'h7f6; 
SIN_ROM[1086] <= 12'h7f6; 
SIN_ROM[1087] <= 12'h7f5; 
SIN_ROM[1088] <= 12'h7f5; 
SIN_ROM[1089] <= 12'h7f5; 
SIN_ROM[1090] <= 12'h7f5; 
SIN_ROM[1091] <= 12'h7f4; 
SIN_ROM[1092] <= 12'h7f4; 
SIN_ROM[1093] <= 12'h7f4; 
SIN_ROM[1094] <= 12'h7f3; 
SIN_ROM[1095] <= 12'h7f3; 
SIN_ROM[1096] <= 12'h7f3; 
SIN_ROM[1097] <= 12'h7f2; 
SIN_ROM[1098] <= 12'h7f2; 
SIN_ROM[1099] <= 12'h7f1; 
SIN_ROM[1100] <= 12'h7f1; 
SIN_ROM[1101] <= 12'h7f1; 
SIN_ROM[1102] <= 12'h7f0; 
SIN_ROM[1103] <= 12'h7f0; 
SIN_ROM[1104] <= 12'h7f0; 
SIN_ROM[1105] <= 12'h7ef; 
SIN_ROM[1106] <= 12'h7ef; 
SIN_ROM[1107] <= 12'h7ee; 
SIN_ROM[1108] <= 12'h7ee; 
SIN_ROM[1109] <= 12'h7ee; 
SIN_ROM[1110] <= 12'h7ed; 
SIN_ROM[1111] <= 12'h7ed; 
SIN_ROM[1112] <= 12'h7ec; 
SIN_ROM[1113] <= 12'h7ec; 
SIN_ROM[1114] <= 12'h7ec; 
SIN_ROM[1115] <= 12'h7eb; 
SIN_ROM[1116] <= 12'h7eb; 
SIN_ROM[1117] <= 12'h7ea; 
SIN_ROM[1118] <= 12'h7ea; 
SIN_ROM[1119] <= 12'h7e9; 
SIN_ROM[1120] <= 12'h7e9; 
SIN_ROM[1121] <= 12'h7e8; 
SIN_ROM[1122] <= 12'h7e8; 
SIN_ROM[1123] <= 12'h7e7; 
SIN_ROM[1124] <= 12'h7e7; 
SIN_ROM[1125] <= 12'h7e6; 
SIN_ROM[1126] <= 12'h7e6; 
SIN_ROM[1127] <= 12'h7e6; 
SIN_ROM[1128] <= 12'h7e5; 
SIN_ROM[1129] <= 12'h7e5; 
SIN_ROM[1130] <= 12'h7e4; 
SIN_ROM[1131] <= 12'h7e3; 
SIN_ROM[1132] <= 12'h7e3; 
SIN_ROM[1133] <= 12'h7e2; 
SIN_ROM[1134] <= 12'h7e2; 
SIN_ROM[1135] <= 12'h7e1; 
SIN_ROM[1136] <= 12'h7e1; 
SIN_ROM[1137] <= 12'h7e0; 
SIN_ROM[1138] <= 12'h7e0; 
SIN_ROM[1139] <= 12'h7df; 
SIN_ROM[1140] <= 12'h7df; 
SIN_ROM[1141] <= 12'h7de; 
SIN_ROM[1142] <= 12'h7de; 
SIN_ROM[1143] <= 12'h7dd; 
SIN_ROM[1144] <= 12'h7dc; 
SIN_ROM[1145] <= 12'h7dc; 
SIN_ROM[1146] <= 12'h7db; 
SIN_ROM[1147] <= 12'h7db; 
SIN_ROM[1148] <= 12'h7da; 
SIN_ROM[1149] <= 12'h7d9; 
SIN_ROM[1150] <= 12'h7d9; 
SIN_ROM[1151] <= 12'h7d8; 
SIN_ROM[1152] <= 12'h7d8; 
SIN_ROM[1153] <= 12'h7d7; 
SIN_ROM[1154] <= 12'h7d6; 
SIN_ROM[1155] <= 12'h7d6; 
SIN_ROM[1156] <= 12'h7d5; 
SIN_ROM[1157] <= 12'h7d5; 
SIN_ROM[1158] <= 12'h7d4; 
SIN_ROM[1159] <= 12'h7d3; 
SIN_ROM[1160] <= 12'h7d3; 
SIN_ROM[1161] <= 12'h7d2; 
SIN_ROM[1162] <= 12'h7d1; 
SIN_ROM[1163] <= 12'h7d1; 
SIN_ROM[1164] <= 12'h7d0; 
SIN_ROM[1165] <= 12'h7cf; 
SIN_ROM[1166] <= 12'h7cf; 
SIN_ROM[1167] <= 12'h7ce; 
SIN_ROM[1168] <= 12'h7cd; 
SIN_ROM[1169] <= 12'h7cd; 
SIN_ROM[1170] <= 12'h7cc; 
SIN_ROM[1171] <= 12'h7cb; 
SIN_ROM[1172] <= 12'h7ca; 
SIN_ROM[1173] <= 12'h7ca; 
SIN_ROM[1174] <= 12'h7c9; 
SIN_ROM[1175] <= 12'h7c8; 
SIN_ROM[1176] <= 12'h7c8; 
SIN_ROM[1177] <= 12'h7c7; 
SIN_ROM[1178] <= 12'h7c6; 
SIN_ROM[1179] <= 12'h7c5; 
SIN_ROM[1180] <= 12'h7c5; 
SIN_ROM[1181] <= 12'h7c4; 
SIN_ROM[1182] <= 12'h7c3; 
SIN_ROM[1183] <= 12'h7c2; 
SIN_ROM[1184] <= 12'h7c2; 
SIN_ROM[1185] <= 12'h7c1; 
SIN_ROM[1186] <= 12'h7c0; 
SIN_ROM[1187] <= 12'h7bf; 
SIN_ROM[1188] <= 12'h7bf; 
SIN_ROM[1189] <= 12'h7be; 
SIN_ROM[1190] <= 12'h7bd; 
SIN_ROM[1191] <= 12'h7bc; 
SIN_ROM[1192] <= 12'h7bb; 
SIN_ROM[1193] <= 12'h7bb; 
SIN_ROM[1194] <= 12'h7ba; 
SIN_ROM[1195] <= 12'h7b9; 
SIN_ROM[1196] <= 12'h7b8; 
SIN_ROM[1197] <= 12'h7b7; 
SIN_ROM[1198] <= 12'h7b7; 
SIN_ROM[1199] <= 12'h7b6; 
SIN_ROM[1200] <= 12'h7b5; 
SIN_ROM[1201] <= 12'h7b4; 
SIN_ROM[1202] <= 12'h7b3; 
SIN_ROM[1203] <= 12'h7b2; 
SIN_ROM[1204] <= 12'h7b1; 
SIN_ROM[1205] <= 12'h7b1; 
SIN_ROM[1206] <= 12'h7b0; 
SIN_ROM[1207] <= 12'h7af; 
SIN_ROM[1208] <= 12'h7ae; 
SIN_ROM[1209] <= 12'h7ad; 
SIN_ROM[1210] <= 12'h7ac; 
SIN_ROM[1211] <= 12'h7ab; 
SIN_ROM[1212] <= 12'h7aa; 
SIN_ROM[1213] <= 12'h7aa; 
SIN_ROM[1214] <= 12'h7a9; 
SIN_ROM[1215] <= 12'h7a8; 
SIN_ROM[1216] <= 12'h7a7; 
SIN_ROM[1217] <= 12'h7a6; 
SIN_ROM[1218] <= 12'h7a5; 
SIN_ROM[1219] <= 12'h7a4; 
SIN_ROM[1220] <= 12'h7a3; 
SIN_ROM[1221] <= 12'h7a2; 
SIN_ROM[1222] <= 12'h7a1; 
SIN_ROM[1223] <= 12'h7a0; 
SIN_ROM[1224] <= 12'h79f; 
SIN_ROM[1225] <= 12'h79e; 
SIN_ROM[1226] <= 12'h79e; 
SIN_ROM[1227] <= 12'h79d; 
SIN_ROM[1228] <= 12'h79c; 
SIN_ROM[1229] <= 12'h79b; 
SIN_ROM[1230] <= 12'h79a; 
SIN_ROM[1231] <= 12'h799; 
SIN_ROM[1232] <= 12'h798; 
SIN_ROM[1233] <= 12'h797; 
SIN_ROM[1234] <= 12'h796; 
SIN_ROM[1235] <= 12'h795; 
SIN_ROM[1236] <= 12'h794; 
SIN_ROM[1237] <= 12'h793; 
SIN_ROM[1238] <= 12'h792; 
SIN_ROM[1239] <= 12'h791; 
SIN_ROM[1240] <= 12'h790; 
SIN_ROM[1241] <= 12'h78f; 
SIN_ROM[1242] <= 12'h78e; 
SIN_ROM[1243] <= 12'h78d; 
SIN_ROM[1244] <= 12'h78c; 
SIN_ROM[1245] <= 12'h78a; 
SIN_ROM[1246] <= 12'h789; 
SIN_ROM[1247] <= 12'h788; 
SIN_ROM[1248] <= 12'h787; 
SIN_ROM[1249] <= 12'h786; 
SIN_ROM[1250] <= 12'h785; 
SIN_ROM[1251] <= 12'h784; 
SIN_ROM[1252] <= 12'h783; 
SIN_ROM[1253] <= 12'h782; 
SIN_ROM[1254] <= 12'h781; 
SIN_ROM[1255] <= 12'h780; 
SIN_ROM[1256] <= 12'h77f; 
SIN_ROM[1257] <= 12'h77e; 
SIN_ROM[1258] <= 12'h77d; 
SIN_ROM[1259] <= 12'h77b; 
SIN_ROM[1260] <= 12'h77a; 
SIN_ROM[1261] <= 12'h779; 
SIN_ROM[1262] <= 12'h778; 
SIN_ROM[1263] <= 12'h777; 
SIN_ROM[1264] <= 12'h776; 
SIN_ROM[1265] <= 12'h775; 
SIN_ROM[1266] <= 12'h774; 
SIN_ROM[1267] <= 12'h772; 
SIN_ROM[1268] <= 12'h771; 
SIN_ROM[1269] <= 12'h770; 
SIN_ROM[1270] <= 12'h76f; 
SIN_ROM[1271] <= 12'h76e; 
SIN_ROM[1272] <= 12'h76d; 
SIN_ROM[1273] <= 12'h76b; 
SIN_ROM[1274] <= 12'h76a; 
SIN_ROM[1275] <= 12'h769; 
SIN_ROM[1276] <= 12'h768; 
SIN_ROM[1277] <= 12'h767; 
SIN_ROM[1278] <= 12'h766; 
SIN_ROM[1279] <= 12'h764; 
SIN_ROM[1280] <= 12'h763; 
SIN_ROM[1281] <= 12'h762; 
SIN_ROM[1282] <= 12'h761; 
SIN_ROM[1283] <= 12'h760; 
SIN_ROM[1284] <= 12'h75e; 
SIN_ROM[1285] <= 12'h75d; 
SIN_ROM[1286] <= 12'h75c; 
SIN_ROM[1287] <= 12'h75b; 
SIN_ROM[1288] <= 12'h759; 
SIN_ROM[1289] <= 12'h758; 
SIN_ROM[1290] <= 12'h757; 
SIN_ROM[1291] <= 12'h756; 
SIN_ROM[1292] <= 12'h754; 
SIN_ROM[1293] <= 12'h753; 
SIN_ROM[1294] <= 12'h752; 
SIN_ROM[1295] <= 12'h751; 
SIN_ROM[1296] <= 12'h74f; 
SIN_ROM[1297] <= 12'h74e; 
SIN_ROM[1298] <= 12'h74d; 
SIN_ROM[1299] <= 12'h74c; 
SIN_ROM[1300] <= 12'h74a; 
SIN_ROM[1301] <= 12'h749; 
SIN_ROM[1302] <= 12'h748; 
SIN_ROM[1303] <= 12'h746; 
SIN_ROM[1304] <= 12'h745; 
SIN_ROM[1305] <= 12'h744; 
SIN_ROM[1306] <= 12'h742; 
SIN_ROM[1307] <= 12'h741; 
SIN_ROM[1308] <= 12'h740; 
SIN_ROM[1309] <= 12'h73e; 
SIN_ROM[1310] <= 12'h73d; 
SIN_ROM[1311] <= 12'h73c; 
SIN_ROM[1312] <= 12'h73a; 
SIN_ROM[1313] <= 12'h739; 
SIN_ROM[1314] <= 12'h738; 
SIN_ROM[1315] <= 12'h736; 
SIN_ROM[1316] <= 12'h735; 
SIN_ROM[1317] <= 12'h734; 
SIN_ROM[1318] <= 12'h732; 
SIN_ROM[1319] <= 12'h731; 
SIN_ROM[1320] <= 12'h730; 
SIN_ROM[1321] <= 12'h72e; 
SIN_ROM[1322] <= 12'h72d; 
SIN_ROM[1323] <= 12'h72b; 
SIN_ROM[1324] <= 12'h72a; 
SIN_ROM[1325] <= 12'h729; 
SIN_ROM[1326] <= 12'h727; 
SIN_ROM[1327] <= 12'h726; 
SIN_ROM[1328] <= 12'h724; 
SIN_ROM[1329] <= 12'h723; 
SIN_ROM[1330] <= 12'h722; 
SIN_ROM[1331] <= 12'h720; 
SIN_ROM[1332] <= 12'h71f; 
SIN_ROM[1333] <= 12'h71d; 
SIN_ROM[1334] <= 12'h71c; 
SIN_ROM[1335] <= 12'h71a; 
SIN_ROM[1336] <= 12'h719; 
SIN_ROM[1337] <= 12'h718; 
SIN_ROM[1338] <= 12'h716; 
SIN_ROM[1339] <= 12'h715; 
SIN_ROM[1340] <= 12'h713; 
SIN_ROM[1341] <= 12'h712; 
SIN_ROM[1342] <= 12'h710; 
SIN_ROM[1343] <= 12'h70f; 
SIN_ROM[1344] <= 12'h70d; 
SIN_ROM[1345] <= 12'h70c; 
SIN_ROM[1346] <= 12'h70a; 
SIN_ROM[1347] <= 12'h709; 
SIN_ROM[1348] <= 12'h707; 
SIN_ROM[1349] <= 12'h706; 
SIN_ROM[1350] <= 12'h704; 
SIN_ROM[1351] <= 12'h703; 
SIN_ROM[1352] <= 12'h701; 
SIN_ROM[1353] <= 12'h700; 
SIN_ROM[1354] <= 12'h6fe; 
SIN_ROM[1355] <= 12'h6fd; 
SIN_ROM[1356] <= 12'h6fb; 
SIN_ROM[1357] <= 12'h6fa; 
SIN_ROM[1358] <= 12'h6f8; 
SIN_ROM[1359] <= 12'h6f7; 
SIN_ROM[1360] <= 12'h6f5; 
SIN_ROM[1361] <= 12'h6f4; 
SIN_ROM[1362] <= 12'h6f2; 
SIN_ROM[1363] <= 12'h6f0; 
SIN_ROM[1364] <= 12'h6ef; 
SIN_ROM[1365] <= 12'h6ed; 
SIN_ROM[1366] <= 12'h6ec; 
SIN_ROM[1367] <= 12'h6ea; 
SIN_ROM[1368] <= 12'h6e9; 
SIN_ROM[1369] <= 12'h6e7; 
SIN_ROM[1370] <= 12'h6e5; 
SIN_ROM[1371] <= 12'h6e4; 
SIN_ROM[1372] <= 12'h6e2; 
SIN_ROM[1373] <= 12'h6e1; 
SIN_ROM[1374] <= 12'h6df; 
SIN_ROM[1375] <= 12'h6dd; 
SIN_ROM[1376] <= 12'h6dc; 
SIN_ROM[1377] <= 12'h6da; 
SIN_ROM[1378] <= 12'h6d9; 
SIN_ROM[1379] <= 12'h6d7; 
SIN_ROM[1380] <= 12'h6d5; 
SIN_ROM[1381] <= 12'h6d4; 
SIN_ROM[1382] <= 12'h6d2; 
SIN_ROM[1383] <= 12'h6d0; 
SIN_ROM[1384] <= 12'h6cf; 
SIN_ROM[1385] <= 12'h6cd; 
SIN_ROM[1386] <= 12'h6cb; 
SIN_ROM[1387] <= 12'h6ca; 
SIN_ROM[1388] <= 12'h6c8; 
SIN_ROM[1389] <= 12'h6c6; 
SIN_ROM[1390] <= 12'h6c5; 
SIN_ROM[1391] <= 12'h6c3; 
SIN_ROM[1392] <= 12'h6c1; 
SIN_ROM[1393] <= 12'h6c0; 
SIN_ROM[1394] <= 12'h6be; 
SIN_ROM[1395] <= 12'h6bc; 
SIN_ROM[1396] <= 12'h6bb; 
SIN_ROM[1397] <= 12'h6b9; 
SIN_ROM[1398] <= 12'h6b7; 
SIN_ROM[1399] <= 12'h6b6; 
SIN_ROM[1400] <= 12'h6b4; 
SIN_ROM[1401] <= 12'h6b2; 
SIN_ROM[1402] <= 12'h6b0; 
SIN_ROM[1403] <= 12'h6af; 
SIN_ROM[1404] <= 12'h6ad; 
SIN_ROM[1405] <= 12'h6ab; 
SIN_ROM[1406] <= 12'h6a9; 
SIN_ROM[1407] <= 12'h6a8; 
SIN_ROM[1408] <= 12'h6a6; 
SIN_ROM[1409] <= 12'h6a4; 
SIN_ROM[1410] <= 12'h6a3; 
SIN_ROM[1411] <= 12'h6a1; 
SIN_ROM[1412] <= 12'h69f; 
SIN_ROM[1413] <= 12'h69d; 
SIN_ROM[1414] <= 12'h69b; 
SIN_ROM[1415] <= 12'h69a; 
SIN_ROM[1416] <= 12'h698; 
SIN_ROM[1417] <= 12'h696; 
SIN_ROM[1418] <= 12'h694; 
SIN_ROM[1419] <= 12'h693; 
SIN_ROM[1420] <= 12'h691; 
SIN_ROM[1421] <= 12'h68f; 
SIN_ROM[1422] <= 12'h68d; 
SIN_ROM[1423] <= 12'h68b; 
SIN_ROM[1424] <= 12'h68a; 
SIN_ROM[1425] <= 12'h688; 
SIN_ROM[1426] <= 12'h686; 
SIN_ROM[1427] <= 12'h684; 
SIN_ROM[1428] <= 12'h682; 
SIN_ROM[1429] <= 12'h681; 
SIN_ROM[1430] <= 12'h67f; 
SIN_ROM[1431] <= 12'h67d; 
SIN_ROM[1432] <= 12'h67b; 
SIN_ROM[1433] <= 12'h679; 
SIN_ROM[1434] <= 12'h677; 
SIN_ROM[1435] <= 12'h675; 
SIN_ROM[1436] <= 12'h674; 
SIN_ROM[1437] <= 12'h672; 
SIN_ROM[1438] <= 12'h670; 
SIN_ROM[1439] <= 12'h66e; 
SIN_ROM[1440] <= 12'h66c; 
SIN_ROM[1441] <= 12'h66a; 
SIN_ROM[1442] <= 12'h668; 
SIN_ROM[1443] <= 12'h667; 
SIN_ROM[1444] <= 12'h665; 
SIN_ROM[1445] <= 12'h663; 
SIN_ROM[1446] <= 12'h661; 
SIN_ROM[1447] <= 12'h65f; 
SIN_ROM[1448] <= 12'h65d; 
SIN_ROM[1449] <= 12'h65b; 
SIN_ROM[1450] <= 12'h659; 
SIN_ROM[1451] <= 12'h657; 
SIN_ROM[1452] <= 12'h655; 
SIN_ROM[1453] <= 12'h654; 
SIN_ROM[1454] <= 12'h652; 
SIN_ROM[1455] <= 12'h650; 
SIN_ROM[1456] <= 12'h64e; 
SIN_ROM[1457] <= 12'h64c; 
SIN_ROM[1458] <= 12'h64a; 
SIN_ROM[1459] <= 12'h648; 
SIN_ROM[1460] <= 12'h646; 
SIN_ROM[1461] <= 12'h644; 
SIN_ROM[1462] <= 12'h642; 
SIN_ROM[1463] <= 12'h640; 
SIN_ROM[1464] <= 12'h63e; 
SIN_ROM[1465] <= 12'h63c; 
SIN_ROM[1466] <= 12'h63a; 
SIN_ROM[1467] <= 12'h638; 
SIN_ROM[1468] <= 12'h636; 
SIN_ROM[1469] <= 12'h634; 
SIN_ROM[1470] <= 12'h632; 
SIN_ROM[1471] <= 12'h630; 
SIN_ROM[1472] <= 12'h62e; 
SIN_ROM[1473] <= 12'h62c; 
SIN_ROM[1474] <= 12'h62a; 
SIN_ROM[1475] <= 12'h628; 
SIN_ROM[1476] <= 12'h626; 
SIN_ROM[1477] <= 12'h624; 
SIN_ROM[1478] <= 12'h622; 
SIN_ROM[1479] <= 12'h620; 
SIN_ROM[1480] <= 12'h61e; 
SIN_ROM[1481] <= 12'h61c; 
SIN_ROM[1482] <= 12'h61a; 
SIN_ROM[1483] <= 12'h618; 
SIN_ROM[1484] <= 12'h616; 
SIN_ROM[1485] <= 12'h614; 
SIN_ROM[1486] <= 12'h612; 
SIN_ROM[1487] <= 12'h610; 
SIN_ROM[1488] <= 12'h60e; 
SIN_ROM[1489] <= 12'h60c; 
SIN_ROM[1490] <= 12'h60a; 
SIN_ROM[1491] <= 12'h608; 
SIN_ROM[1492] <= 12'h606; 
SIN_ROM[1493] <= 12'h604; 
SIN_ROM[1494] <= 12'h602; 
SIN_ROM[1495] <= 12'h600; 
SIN_ROM[1496] <= 12'h5fd; 
SIN_ROM[1497] <= 12'h5fb; 
SIN_ROM[1498] <= 12'h5f9; 
SIN_ROM[1499] <= 12'h5f7; 
SIN_ROM[1500] <= 12'h5f5; 
SIN_ROM[1501] <= 12'h5f3; 
SIN_ROM[1502] <= 12'h5f1; 
SIN_ROM[1503] <= 12'h5ef; 
SIN_ROM[1504] <= 12'h5ed; 
SIN_ROM[1505] <= 12'h5eb; 
SIN_ROM[1506] <= 12'h5e9; 
SIN_ROM[1507] <= 12'h5e6; 
SIN_ROM[1508] <= 12'h5e4; 
SIN_ROM[1509] <= 12'h5e2; 
SIN_ROM[1510] <= 12'h5e0; 
SIN_ROM[1511] <= 12'h5de; 
SIN_ROM[1512] <= 12'h5dc; 
SIN_ROM[1513] <= 12'h5da; 
SIN_ROM[1514] <= 12'h5d7; 
SIN_ROM[1515] <= 12'h5d5; 
SIN_ROM[1516] <= 12'h5d3; 
SIN_ROM[1517] <= 12'h5d1; 
SIN_ROM[1518] <= 12'h5cf; 
SIN_ROM[1519] <= 12'h5cd; 
SIN_ROM[1520] <= 12'h5cb; 
SIN_ROM[1521] <= 12'h5c8; 
SIN_ROM[1522] <= 12'h5c6; 
SIN_ROM[1523] <= 12'h5c4; 
SIN_ROM[1524] <= 12'h5c2; 
SIN_ROM[1525] <= 12'h5c0; 
SIN_ROM[1526] <= 12'h5bd; 
SIN_ROM[1527] <= 12'h5bb; 
SIN_ROM[1528] <= 12'h5b9; 
SIN_ROM[1529] <= 12'h5b7; 
SIN_ROM[1530] <= 12'h5b5; 
SIN_ROM[1531] <= 12'h5b3; 
SIN_ROM[1532] <= 12'h5b0; 
SIN_ROM[1533] <= 12'h5ae; 
SIN_ROM[1534] <= 12'h5ac; 
SIN_ROM[1535] <= 12'h5aa; 
SIN_ROM[1536] <= 12'h5a7; 
SIN_ROM[1537] <= 12'h5a5; 
SIN_ROM[1538] <= 12'h5a3; 
SIN_ROM[1539] <= 12'h5a1; 
SIN_ROM[1540] <= 12'h59f; 
SIN_ROM[1541] <= 12'h59c; 
SIN_ROM[1542] <= 12'h59a; 
SIN_ROM[1543] <= 12'h598; 
SIN_ROM[1544] <= 12'h596; 
SIN_ROM[1545] <= 12'h593; 
SIN_ROM[1546] <= 12'h591; 
SIN_ROM[1547] <= 12'h58f; 
SIN_ROM[1548] <= 12'h58d; 
SIN_ROM[1549] <= 12'h58a; 
SIN_ROM[1550] <= 12'h588; 
SIN_ROM[1551] <= 12'h586; 
SIN_ROM[1552] <= 12'h583; 
SIN_ROM[1553] <= 12'h581; 
SIN_ROM[1554] <= 12'h57f; 
SIN_ROM[1555] <= 12'h57d; 
SIN_ROM[1556] <= 12'h57a; 
SIN_ROM[1557] <= 12'h578; 
SIN_ROM[1558] <= 12'h576; 
SIN_ROM[1559] <= 12'h573; 
SIN_ROM[1560] <= 12'h571; 
SIN_ROM[1561] <= 12'h56f; 
SIN_ROM[1562] <= 12'h56d; 
SIN_ROM[1563] <= 12'h56a; 
SIN_ROM[1564] <= 12'h568; 
SIN_ROM[1565] <= 12'h566; 
SIN_ROM[1566] <= 12'h563; 
SIN_ROM[1567] <= 12'h561; 
SIN_ROM[1568] <= 12'h55f; 
SIN_ROM[1569] <= 12'h55c; 
SIN_ROM[1570] <= 12'h55a; 
SIN_ROM[1571] <= 12'h558; 
SIN_ROM[1572] <= 12'h555; 
SIN_ROM[1573] <= 12'h553; 
SIN_ROM[1574] <= 12'h551; 
SIN_ROM[1575] <= 12'h54e; 
SIN_ROM[1576] <= 12'h54c; 
SIN_ROM[1577] <= 12'h54a; 
SIN_ROM[1578] <= 12'h547; 
SIN_ROM[1579] <= 12'h545; 
SIN_ROM[1580] <= 12'h543; 
SIN_ROM[1581] <= 12'h540; 
SIN_ROM[1582] <= 12'h53e; 
SIN_ROM[1583] <= 12'h53b; 
SIN_ROM[1584] <= 12'h539; 
SIN_ROM[1585] <= 12'h537; 
SIN_ROM[1586] <= 12'h534; 
SIN_ROM[1587] <= 12'h532; 
SIN_ROM[1588] <= 12'h530; 
SIN_ROM[1589] <= 12'h52d; 
SIN_ROM[1590] <= 12'h52b; 
SIN_ROM[1591] <= 12'h528; 
SIN_ROM[1592] <= 12'h526; 
SIN_ROM[1593] <= 12'h524; 
SIN_ROM[1594] <= 12'h521; 
SIN_ROM[1595] <= 12'h51f; 
SIN_ROM[1596] <= 12'h51c; 
SIN_ROM[1597] <= 12'h51a; 
SIN_ROM[1598] <= 12'h517; 
SIN_ROM[1599] <= 12'h515; 
SIN_ROM[1600] <= 12'h513; 
SIN_ROM[1601] <= 12'h510; 
SIN_ROM[1602] <= 12'h50e; 
SIN_ROM[1603] <= 12'h50b; 
SIN_ROM[1604] <= 12'h509; 
SIN_ROM[1605] <= 12'h506; 
SIN_ROM[1606] <= 12'h504; 
SIN_ROM[1607] <= 12'h502; 
SIN_ROM[1608] <= 12'h4ff; 
SIN_ROM[1609] <= 12'h4fd; 
SIN_ROM[1610] <= 12'h4fa; 
SIN_ROM[1611] <= 12'h4f8; 
SIN_ROM[1612] <= 12'h4f5; 
SIN_ROM[1613] <= 12'h4f3; 
SIN_ROM[1614] <= 12'h4f0; 
SIN_ROM[1615] <= 12'h4ee; 
SIN_ROM[1616] <= 12'h4eb; 
SIN_ROM[1617] <= 12'h4e9; 
SIN_ROM[1618] <= 12'h4e6; 
SIN_ROM[1619] <= 12'h4e4; 
SIN_ROM[1620] <= 12'h4e1; 
SIN_ROM[1621] <= 12'h4df; 
SIN_ROM[1622] <= 12'h4dc; 
SIN_ROM[1623] <= 12'h4da; 
SIN_ROM[1624] <= 12'h4d7; 
SIN_ROM[1625] <= 12'h4d5; 
SIN_ROM[1626] <= 12'h4d2; 
SIN_ROM[1627] <= 12'h4d0; 
SIN_ROM[1628] <= 12'h4cd; 
SIN_ROM[1629] <= 12'h4cb; 
SIN_ROM[1630] <= 12'h4c8; 
SIN_ROM[1631] <= 12'h4c6; 
SIN_ROM[1632] <= 12'h4c3; 
SIN_ROM[1633] <= 12'h4c1; 
SIN_ROM[1634] <= 12'h4be; 
SIN_ROM[1635] <= 12'h4bc; 
SIN_ROM[1636] <= 12'h4b9; 
SIN_ROM[1637] <= 12'h4b7; 
SIN_ROM[1638] <= 12'h4b4; 
SIN_ROM[1639] <= 12'h4b2; 
SIN_ROM[1640] <= 12'h4af; 
SIN_ROM[1641] <= 12'h4ad; 
SIN_ROM[1642] <= 12'h4aa; 
SIN_ROM[1643] <= 12'h4a7; 
SIN_ROM[1644] <= 12'h4a5; 
SIN_ROM[1645] <= 12'h4a2; 
SIN_ROM[1646] <= 12'h4a0; 
SIN_ROM[1647] <= 12'h49d; 
SIN_ROM[1648] <= 12'h49b; 
SIN_ROM[1649] <= 12'h498; 
SIN_ROM[1650] <= 12'h496; 
SIN_ROM[1651] <= 12'h493; 
SIN_ROM[1652] <= 12'h490; 
SIN_ROM[1653] <= 12'h48e; 
SIN_ROM[1654] <= 12'h48b; 
SIN_ROM[1655] <= 12'h489; 
SIN_ROM[1656] <= 12'h486; 
SIN_ROM[1657] <= 12'h483; 
SIN_ROM[1658] <= 12'h481; 
SIN_ROM[1659] <= 12'h47e; 
SIN_ROM[1660] <= 12'h47c; 
SIN_ROM[1661] <= 12'h479; 
SIN_ROM[1662] <= 12'h476; 
SIN_ROM[1663] <= 12'h474; 
SIN_ROM[1664] <= 12'h471; 
SIN_ROM[1665] <= 12'h46f; 
SIN_ROM[1666] <= 12'h46c; 
SIN_ROM[1667] <= 12'h469; 
SIN_ROM[1668] <= 12'h467; 
SIN_ROM[1669] <= 12'h464; 
SIN_ROM[1670] <= 12'h462; 
SIN_ROM[1671] <= 12'h45f; 
SIN_ROM[1672] <= 12'h45c; 
SIN_ROM[1673] <= 12'h45a; 
SIN_ROM[1674] <= 12'h457; 
SIN_ROM[1675] <= 12'h454; 
SIN_ROM[1676] <= 12'h452; 
SIN_ROM[1677] <= 12'h44f; 
SIN_ROM[1678] <= 12'h44c; 
SIN_ROM[1679] <= 12'h44a; 
SIN_ROM[1680] <= 12'h447; 
SIN_ROM[1681] <= 12'h444; 
SIN_ROM[1682] <= 12'h442; 
SIN_ROM[1683] <= 12'h43f; 
SIN_ROM[1684] <= 12'h43d; 
SIN_ROM[1685] <= 12'h43a; 
SIN_ROM[1686] <= 12'h437; 
SIN_ROM[1687] <= 12'h435; 
SIN_ROM[1688] <= 12'h432; 
SIN_ROM[1689] <= 12'h42f; 
SIN_ROM[1690] <= 12'h42c; 
SIN_ROM[1691] <= 12'h42a; 
SIN_ROM[1692] <= 12'h427; 
SIN_ROM[1693] <= 12'h424; 
SIN_ROM[1694] <= 12'h422; 
SIN_ROM[1695] <= 12'h41f; 
SIN_ROM[1696] <= 12'h41c; 
SIN_ROM[1697] <= 12'h41a; 
SIN_ROM[1698] <= 12'h417; 
SIN_ROM[1699] <= 12'h414; 
SIN_ROM[1700] <= 12'h412; 
SIN_ROM[1701] <= 12'h40f; 
SIN_ROM[1702] <= 12'h40c; 
SIN_ROM[1703] <= 12'h409; 
SIN_ROM[1704] <= 12'h407; 
SIN_ROM[1705] <= 12'h404; 
SIN_ROM[1706] <= 12'h401; 
SIN_ROM[1707] <= 12'h3ff; 
SIN_ROM[1708] <= 12'h3fc; 
SIN_ROM[1709] <= 12'h3f9; 
SIN_ROM[1710] <= 12'h3f6; 
SIN_ROM[1711] <= 12'h3f4; 
SIN_ROM[1712] <= 12'h3f1; 
SIN_ROM[1713] <= 12'h3ee; 
SIN_ROM[1714] <= 12'h3eb; 
SIN_ROM[1715] <= 12'h3e9; 
SIN_ROM[1716] <= 12'h3e6; 
SIN_ROM[1717] <= 12'h3e3; 
SIN_ROM[1718] <= 12'h3e1; 
SIN_ROM[1719] <= 12'h3de; 
SIN_ROM[1720] <= 12'h3db; 
SIN_ROM[1721] <= 12'h3d8; 
SIN_ROM[1722] <= 12'h3d6; 
SIN_ROM[1723] <= 12'h3d3; 
SIN_ROM[1724] <= 12'h3d0; 
SIN_ROM[1725] <= 12'h3cd; 
SIN_ROM[1726] <= 12'h3ca; 
SIN_ROM[1727] <= 12'h3c8; 
SIN_ROM[1728] <= 12'h3c5; 
SIN_ROM[1729] <= 12'h3c2; 
SIN_ROM[1730] <= 12'h3bf; 
SIN_ROM[1731] <= 12'h3bd; 
SIN_ROM[1732] <= 12'h3ba; 
SIN_ROM[1733] <= 12'h3b7; 
SIN_ROM[1734] <= 12'h3b4; 
SIN_ROM[1735] <= 12'h3b2; 
SIN_ROM[1736] <= 12'h3af; 
SIN_ROM[1737] <= 12'h3ac; 
SIN_ROM[1738] <= 12'h3a9; 
SIN_ROM[1739] <= 12'h3a6; 
SIN_ROM[1740] <= 12'h3a4; 
SIN_ROM[1741] <= 12'h3a1; 
SIN_ROM[1742] <= 12'h39e; 
SIN_ROM[1743] <= 12'h39b; 
SIN_ROM[1744] <= 12'h398; 
SIN_ROM[1745] <= 12'h396; 
SIN_ROM[1746] <= 12'h393; 
SIN_ROM[1747] <= 12'h390; 
SIN_ROM[1748] <= 12'h38d; 
SIN_ROM[1749] <= 12'h38a; 
SIN_ROM[1750] <= 12'h387; 
SIN_ROM[1751] <= 12'h385; 
SIN_ROM[1752] <= 12'h382; 
SIN_ROM[1753] <= 12'h37f; 
SIN_ROM[1754] <= 12'h37c; 
SIN_ROM[1755] <= 12'h379; 
SIN_ROM[1756] <= 12'h377; 
SIN_ROM[1757] <= 12'h374; 
SIN_ROM[1758] <= 12'h371; 
SIN_ROM[1759] <= 12'h36e; 
SIN_ROM[1760] <= 12'h36b; 
SIN_ROM[1761] <= 12'h368; 
SIN_ROM[1762] <= 12'h366; 
SIN_ROM[1763] <= 12'h363; 
SIN_ROM[1764] <= 12'h360; 
SIN_ROM[1765] <= 12'h35d; 
SIN_ROM[1766] <= 12'h35a; 
SIN_ROM[1767] <= 12'h357; 
SIN_ROM[1768] <= 12'h354; 
SIN_ROM[1769] <= 12'h352; 
SIN_ROM[1770] <= 12'h34f; 
SIN_ROM[1771] <= 12'h34c; 
SIN_ROM[1772] <= 12'h349; 
SIN_ROM[1773] <= 12'h346; 
SIN_ROM[1774] <= 12'h343; 
SIN_ROM[1775] <= 12'h340; 
SIN_ROM[1776] <= 12'h33e; 
SIN_ROM[1777] <= 12'h33b; 
SIN_ROM[1778] <= 12'h338; 
SIN_ROM[1779] <= 12'h335; 
SIN_ROM[1780] <= 12'h332; 
SIN_ROM[1781] <= 12'h32f; 
SIN_ROM[1782] <= 12'h32c; 
SIN_ROM[1783] <= 12'h329; 
SIN_ROM[1784] <= 12'h327; 
SIN_ROM[1785] <= 12'h324; 
SIN_ROM[1786] <= 12'h321; 
SIN_ROM[1787] <= 12'h31e; 
SIN_ROM[1788] <= 12'h31b; 
SIN_ROM[1789] <= 12'h318; 
SIN_ROM[1790] <= 12'h315; 
SIN_ROM[1791] <= 12'h312; 
SIN_ROM[1792] <= 12'h30f; 
SIN_ROM[1793] <= 12'h30c; 
SIN_ROM[1794] <= 12'h30a; 
SIN_ROM[1795] <= 12'h307; 
SIN_ROM[1796] <= 12'h304; 
SIN_ROM[1797] <= 12'h301; 
SIN_ROM[1798] <= 12'h2fe; 
SIN_ROM[1799] <= 12'h2fb; 
SIN_ROM[1800] <= 12'h2f8; 
SIN_ROM[1801] <= 12'h2f5; 
SIN_ROM[1802] <= 12'h2f2; 
SIN_ROM[1803] <= 12'h2ef; 
SIN_ROM[1804] <= 12'h2ec; 
SIN_ROM[1805] <= 12'h2e9; 
SIN_ROM[1806] <= 12'h2e7; 
SIN_ROM[1807] <= 12'h2e4; 
SIN_ROM[1808] <= 12'h2e1; 
SIN_ROM[1809] <= 12'h2de; 
SIN_ROM[1810] <= 12'h2db; 
SIN_ROM[1811] <= 12'h2d8; 
SIN_ROM[1812] <= 12'h2d5; 
SIN_ROM[1813] <= 12'h2d2; 
SIN_ROM[1814] <= 12'h2cf; 
SIN_ROM[1815] <= 12'h2cc; 
SIN_ROM[1816] <= 12'h2c9; 
SIN_ROM[1817] <= 12'h2c6; 
SIN_ROM[1818] <= 12'h2c3; 
SIN_ROM[1819] <= 12'h2c0; 
SIN_ROM[1820] <= 12'h2bd; 
SIN_ROM[1821] <= 12'h2ba; 
SIN_ROM[1822] <= 12'h2b8; 
SIN_ROM[1823] <= 12'h2b5; 
SIN_ROM[1824] <= 12'h2b2; 
SIN_ROM[1825] <= 12'h2af; 
SIN_ROM[1826] <= 12'h2ac; 
SIN_ROM[1827] <= 12'h2a9; 
SIN_ROM[1828] <= 12'h2a6; 
SIN_ROM[1829] <= 12'h2a3; 
SIN_ROM[1830] <= 12'h2a0; 
SIN_ROM[1831] <= 12'h29d; 
SIN_ROM[1832] <= 12'h29a; 
SIN_ROM[1833] <= 12'h297; 
SIN_ROM[1834] <= 12'h294; 
SIN_ROM[1835] <= 12'h291; 
SIN_ROM[1836] <= 12'h28e; 
SIN_ROM[1837] <= 12'h28b; 
SIN_ROM[1838] <= 12'h288; 
SIN_ROM[1839] <= 12'h285; 
SIN_ROM[1840] <= 12'h282; 
SIN_ROM[1841] <= 12'h27f; 
SIN_ROM[1842] <= 12'h27c; 
SIN_ROM[1843] <= 12'h279; 
SIN_ROM[1844] <= 12'h276; 
SIN_ROM[1845] <= 12'h273; 
SIN_ROM[1846] <= 12'h270; 
SIN_ROM[1847] <= 12'h26d; 
SIN_ROM[1848] <= 12'h26a; 
SIN_ROM[1849] <= 12'h267; 
SIN_ROM[1850] <= 12'h264; 
SIN_ROM[1851] <= 12'h261; 
SIN_ROM[1852] <= 12'h25e; 
SIN_ROM[1853] <= 12'h25b; 
SIN_ROM[1854] <= 12'h258; 
SIN_ROM[1855] <= 12'h255; 
SIN_ROM[1856] <= 12'h252; 
SIN_ROM[1857] <= 12'h24f; 
SIN_ROM[1858] <= 12'h24c; 
SIN_ROM[1859] <= 12'h249; 
SIN_ROM[1860] <= 12'h246; 
SIN_ROM[1861] <= 12'h243; 
SIN_ROM[1862] <= 12'h240; 
SIN_ROM[1863] <= 12'h23d; 
SIN_ROM[1864] <= 12'h23a; 
SIN_ROM[1865] <= 12'h237; 
SIN_ROM[1866] <= 12'h234; 
SIN_ROM[1867] <= 12'h231; 
SIN_ROM[1868] <= 12'h22e; 
SIN_ROM[1869] <= 12'h22b; 
SIN_ROM[1870] <= 12'h228; 
SIN_ROM[1871] <= 12'h225; 
SIN_ROM[1872] <= 12'h222; 
SIN_ROM[1873] <= 12'h21f; 
SIN_ROM[1874] <= 12'h21c; 
SIN_ROM[1875] <= 12'h219; 
SIN_ROM[1876] <= 12'h216; 
SIN_ROM[1877] <= 12'h213; 
SIN_ROM[1878] <= 12'h210; 
SIN_ROM[1879] <= 12'h20d; 
SIN_ROM[1880] <= 12'h20a; 
SIN_ROM[1881] <= 12'h207; 
SIN_ROM[1882] <= 12'h204; 
SIN_ROM[1883] <= 12'h201; 
SIN_ROM[1884] <= 12'h1fe; 
SIN_ROM[1885] <= 12'h1fb; 
SIN_ROM[1886] <= 12'h1f7; 
SIN_ROM[1887] <= 12'h1f4; 
SIN_ROM[1888] <= 12'h1f1; 
SIN_ROM[1889] <= 12'h1ee; 
SIN_ROM[1890] <= 12'h1eb; 
SIN_ROM[1891] <= 12'h1e8; 
SIN_ROM[1892] <= 12'h1e5; 
SIN_ROM[1893] <= 12'h1e2; 
SIN_ROM[1894] <= 12'h1df; 
SIN_ROM[1895] <= 12'h1dc; 
SIN_ROM[1896] <= 12'h1d9; 
SIN_ROM[1897] <= 12'h1d6; 
SIN_ROM[1898] <= 12'h1d3; 
SIN_ROM[1899] <= 12'h1d0; 
SIN_ROM[1900] <= 12'h1cd; 
SIN_ROM[1901] <= 12'h1ca; 
SIN_ROM[1902] <= 12'h1c7; 
SIN_ROM[1903] <= 12'h1c4; 
SIN_ROM[1904] <= 12'h1c1; 
SIN_ROM[1905] <= 12'h1bd; 
SIN_ROM[1906] <= 12'h1ba; 
SIN_ROM[1907] <= 12'h1b7; 
SIN_ROM[1908] <= 12'h1b4; 
SIN_ROM[1909] <= 12'h1b1; 
SIN_ROM[1910] <= 12'h1ae; 
SIN_ROM[1911] <= 12'h1ab; 
SIN_ROM[1912] <= 12'h1a8; 
SIN_ROM[1913] <= 12'h1a5; 
SIN_ROM[1914] <= 12'h1a2; 
SIN_ROM[1915] <= 12'h19f; 
SIN_ROM[1916] <= 12'h19c; 
SIN_ROM[1917] <= 12'h199; 
SIN_ROM[1918] <= 12'h196; 
SIN_ROM[1919] <= 12'h192; 
SIN_ROM[1920] <= 12'h18f; 
SIN_ROM[1921] <= 12'h18c; 
SIN_ROM[1922] <= 12'h189; 
SIN_ROM[1923] <= 12'h186; 
SIN_ROM[1924] <= 12'h183; 
SIN_ROM[1925] <= 12'h180; 
SIN_ROM[1926] <= 12'h17d; 
SIN_ROM[1927] <= 12'h17a; 
SIN_ROM[1928] <= 12'h177; 
SIN_ROM[1929] <= 12'h174; 
SIN_ROM[1930] <= 12'h171; 
SIN_ROM[1931] <= 12'h16d; 
SIN_ROM[1932] <= 12'h16a; 
SIN_ROM[1933] <= 12'h167; 
SIN_ROM[1934] <= 12'h164; 
SIN_ROM[1935] <= 12'h161; 
SIN_ROM[1936] <= 12'h15e; 
SIN_ROM[1937] <= 12'h15b; 
SIN_ROM[1938] <= 12'h158; 
SIN_ROM[1939] <= 12'h155; 
SIN_ROM[1940] <= 12'h152; 
SIN_ROM[1941] <= 12'h14e; 
SIN_ROM[1942] <= 12'h14b; 
SIN_ROM[1943] <= 12'h148; 
SIN_ROM[1944] <= 12'h145; 
SIN_ROM[1945] <= 12'h142; 
SIN_ROM[1946] <= 12'h13f; 
SIN_ROM[1947] <= 12'h13c; 
SIN_ROM[1948] <= 12'h139; 
SIN_ROM[1949] <= 12'h136; 
SIN_ROM[1950] <= 12'h133; 
SIN_ROM[1951] <= 12'h12f; 
SIN_ROM[1952] <= 12'h12c; 
SIN_ROM[1953] <= 12'h129; 
SIN_ROM[1954] <= 12'h126; 
SIN_ROM[1955] <= 12'h123; 
SIN_ROM[1956] <= 12'h120; 
SIN_ROM[1957] <= 12'h11d; 
SIN_ROM[1958] <= 12'h11a; 
SIN_ROM[1959] <= 12'h117; 
SIN_ROM[1960] <= 12'h113; 
SIN_ROM[1961] <= 12'h110; 
SIN_ROM[1962] <= 12'h10d; 
SIN_ROM[1963] <= 12'h10a; 
SIN_ROM[1964] <= 12'h107; 
SIN_ROM[1965] <= 12'h104; 
SIN_ROM[1966] <= 12'h101; 
SIN_ROM[1967] <= 12'h0fe; 
SIN_ROM[1968] <= 12'h0fb; 
SIN_ROM[1969] <= 12'h0f7; 
SIN_ROM[1970] <= 12'h0f4; 
SIN_ROM[1971] <= 12'h0f1; 
SIN_ROM[1972] <= 12'h0ee; 
SIN_ROM[1973] <= 12'h0eb; 
SIN_ROM[1974] <= 12'h0e8; 
SIN_ROM[1975] <= 12'h0e5; 
SIN_ROM[1976] <= 12'h0e2; 
SIN_ROM[1977] <= 12'h0df; 
SIN_ROM[1978] <= 12'h0db; 
SIN_ROM[1979] <= 12'h0d8; 
SIN_ROM[1980] <= 12'h0d5; 
SIN_ROM[1981] <= 12'h0d2; 
SIN_ROM[1982] <= 12'h0cf; 
SIN_ROM[1983] <= 12'h0cc; 
SIN_ROM[1984] <= 12'h0c9; 
SIN_ROM[1985] <= 12'h0c6; 
SIN_ROM[1986] <= 12'h0c2; 
SIN_ROM[1987] <= 12'h0bf; 
SIN_ROM[1988] <= 12'h0bc; 
SIN_ROM[1989] <= 12'h0b9; 
SIN_ROM[1990] <= 12'h0b6; 
SIN_ROM[1991] <= 12'h0b3; 
SIN_ROM[1992] <= 12'h0b0; 
SIN_ROM[1993] <= 12'h0ac; 
SIN_ROM[1994] <= 12'h0a9; 
SIN_ROM[1995] <= 12'h0a6; 
SIN_ROM[1996] <= 12'h0a3; 
SIN_ROM[1997] <= 12'h0a0; 
SIN_ROM[1998] <= 12'h09d; 
SIN_ROM[1999] <= 12'h09a; 
SIN_ROM[2000] <= 12'h097; 
SIN_ROM[2001] <= 12'h093; 
SIN_ROM[2002] <= 12'h090; 
SIN_ROM[2003] <= 12'h08d; 
SIN_ROM[2004] <= 12'h08a; 
SIN_ROM[2005] <= 12'h087; 
SIN_ROM[2006] <= 12'h084; 
SIN_ROM[2007] <= 12'h081; 
SIN_ROM[2008] <= 12'h07e; 
SIN_ROM[2009] <= 12'h07a; 
SIN_ROM[2010] <= 12'h077; 
SIN_ROM[2011] <= 12'h074; 
SIN_ROM[2012] <= 12'h071; 
SIN_ROM[2013] <= 12'h06e; 
SIN_ROM[2014] <= 12'h06b; 
SIN_ROM[2015] <= 12'h068; 
SIN_ROM[2016] <= 12'h064; 
SIN_ROM[2017] <= 12'h061; 
SIN_ROM[2018] <= 12'h05e; 
SIN_ROM[2019] <= 12'h05b; 
SIN_ROM[2020] <= 12'h058; 
SIN_ROM[2021] <= 12'h055; 
SIN_ROM[2022] <= 12'h052; 
SIN_ROM[2023] <= 12'h04e; 
SIN_ROM[2024] <= 12'h04b; 
SIN_ROM[2025] <= 12'h048; 
SIN_ROM[2026] <= 12'h045; 
SIN_ROM[2027] <= 12'h042; 
SIN_ROM[2028] <= 12'h03f; 
SIN_ROM[2029] <= 12'h03c; 
SIN_ROM[2030] <= 12'h039; 
SIN_ROM[2031] <= 12'h035; 
SIN_ROM[2032] <= 12'h032; 
SIN_ROM[2033] <= 12'h02f; 
SIN_ROM[2034] <= 12'h02c; 
SIN_ROM[2035] <= 12'h029; 
SIN_ROM[2036] <= 12'h026; 
SIN_ROM[2037] <= 12'h023; 
SIN_ROM[2038] <= 12'h01f; 
SIN_ROM[2039] <= 12'h01c; 
SIN_ROM[2040] <= 12'h019; 
SIN_ROM[2041] <= 12'h016; 
SIN_ROM[2042] <= 12'h013; 
SIN_ROM[2043] <= 12'h010; 
SIN_ROM[2044] <= 12'h00d; 
SIN_ROM[2045] <= 12'h009; 
SIN_ROM[2046] <= 12'h006; 
SIN_ROM[2047] <= 12'h003; 
SIN_ROM[2048] <= 12'h000; 
SIN_ROM[2049] <= 12'hffd; 
SIN_ROM[2050] <= 12'hffa; 
SIN_ROM[2051] <= 12'hff7; 
SIN_ROM[2052] <= 12'hff3; 
SIN_ROM[2053] <= 12'hff0; 
SIN_ROM[2054] <= 12'hfed; 
SIN_ROM[2055] <= 12'hfea; 
SIN_ROM[2056] <= 12'hfe7; 
SIN_ROM[2057] <= 12'hfe4; 
SIN_ROM[2058] <= 12'hfe1; 
SIN_ROM[2059] <= 12'hfdd; 
SIN_ROM[2060] <= 12'hfda; 
SIN_ROM[2061] <= 12'hfd7; 
SIN_ROM[2062] <= 12'hfd4; 
SIN_ROM[2063] <= 12'hfd1; 
SIN_ROM[2064] <= 12'hfce; 
SIN_ROM[2065] <= 12'hfcb; 
SIN_ROM[2066] <= 12'hfc7; 
SIN_ROM[2067] <= 12'hfc4; 
SIN_ROM[2068] <= 12'hfc1; 
SIN_ROM[2069] <= 12'hfbe; 
SIN_ROM[2070] <= 12'hfbb; 
SIN_ROM[2071] <= 12'hfb8; 
SIN_ROM[2072] <= 12'hfb5; 
SIN_ROM[2073] <= 12'hfb2; 
SIN_ROM[2074] <= 12'hfae; 
SIN_ROM[2075] <= 12'hfab; 
SIN_ROM[2076] <= 12'hfa8; 
SIN_ROM[2077] <= 12'hfa5; 
SIN_ROM[2078] <= 12'hfa2; 
SIN_ROM[2079] <= 12'hf9f; 
SIN_ROM[2080] <= 12'hf9c; 
SIN_ROM[2081] <= 12'hf98; 
SIN_ROM[2082] <= 12'hf95; 
SIN_ROM[2083] <= 12'hf92; 
SIN_ROM[2084] <= 12'hf8f; 
SIN_ROM[2085] <= 12'hf8c; 
SIN_ROM[2086] <= 12'hf89; 
SIN_ROM[2087] <= 12'hf86; 
SIN_ROM[2088] <= 12'hf82; 
SIN_ROM[2089] <= 12'hf7f; 
SIN_ROM[2090] <= 12'hf7c; 
SIN_ROM[2091] <= 12'hf79; 
SIN_ROM[2092] <= 12'hf76; 
SIN_ROM[2093] <= 12'hf73; 
SIN_ROM[2094] <= 12'hf70; 
SIN_ROM[2095] <= 12'hf6d; 
SIN_ROM[2096] <= 12'hf69; 
SIN_ROM[2097] <= 12'hf66; 
SIN_ROM[2098] <= 12'hf63; 
SIN_ROM[2099] <= 12'hf60; 
SIN_ROM[2100] <= 12'hf5d; 
SIN_ROM[2101] <= 12'hf5a; 
SIN_ROM[2102] <= 12'hf57; 
SIN_ROM[2103] <= 12'hf54; 
SIN_ROM[2104] <= 12'hf50; 
SIN_ROM[2105] <= 12'hf4d; 
SIN_ROM[2106] <= 12'hf4a; 
SIN_ROM[2107] <= 12'hf47; 
SIN_ROM[2108] <= 12'hf44; 
SIN_ROM[2109] <= 12'hf41; 
SIN_ROM[2110] <= 12'hf3e; 
SIN_ROM[2111] <= 12'hf3a; 
SIN_ROM[2112] <= 12'hf37; 
SIN_ROM[2113] <= 12'hf34; 
SIN_ROM[2114] <= 12'hf31; 
SIN_ROM[2115] <= 12'hf2e; 
SIN_ROM[2116] <= 12'hf2b; 
SIN_ROM[2117] <= 12'hf28; 
SIN_ROM[2118] <= 12'hf25; 
SIN_ROM[2119] <= 12'hf21; 
SIN_ROM[2120] <= 12'hf1e; 
SIN_ROM[2121] <= 12'hf1b; 
SIN_ROM[2122] <= 12'hf18; 
SIN_ROM[2123] <= 12'hf15; 
SIN_ROM[2124] <= 12'hf12; 
SIN_ROM[2125] <= 12'hf0f; 
SIN_ROM[2126] <= 12'hf0c; 
SIN_ROM[2127] <= 12'hf09; 
SIN_ROM[2128] <= 12'hf05; 
SIN_ROM[2129] <= 12'hf02; 
SIN_ROM[2130] <= 12'heff; 
SIN_ROM[2131] <= 12'hefc; 
SIN_ROM[2132] <= 12'hef9; 
SIN_ROM[2133] <= 12'hef6; 
SIN_ROM[2134] <= 12'hef3; 
SIN_ROM[2135] <= 12'hef0; 
SIN_ROM[2136] <= 12'heed; 
SIN_ROM[2137] <= 12'hee9; 
SIN_ROM[2138] <= 12'hee6; 
SIN_ROM[2139] <= 12'hee3; 
SIN_ROM[2140] <= 12'hee0; 
SIN_ROM[2141] <= 12'hedd; 
SIN_ROM[2142] <= 12'heda; 
SIN_ROM[2143] <= 12'hed7; 
SIN_ROM[2144] <= 12'hed4; 
SIN_ROM[2145] <= 12'hed1; 
SIN_ROM[2146] <= 12'hecd; 
SIN_ROM[2147] <= 12'heca; 
SIN_ROM[2148] <= 12'hec7; 
SIN_ROM[2149] <= 12'hec4; 
SIN_ROM[2150] <= 12'hec1; 
SIN_ROM[2151] <= 12'hebe; 
SIN_ROM[2152] <= 12'hebb; 
SIN_ROM[2153] <= 12'heb8; 
SIN_ROM[2154] <= 12'heb5; 
SIN_ROM[2155] <= 12'heb2; 
SIN_ROM[2156] <= 12'heae; 
SIN_ROM[2157] <= 12'heab; 
SIN_ROM[2158] <= 12'hea8; 
SIN_ROM[2159] <= 12'hea5; 
SIN_ROM[2160] <= 12'hea2; 
SIN_ROM[2161] <= 12'he9f; 
SIN_ROM[2162] <= 12'he9c; 
SIN_ROM[2163] <= 12'he99; 
SIN_ROM[2164] <= 12'he96; 
SIN_ROM[2165] <= 12'he93; 
SIN_ROM[2166] <= 12'he8f; 
SIN_ROM[2167] <= 12'he8c; 
SIN_ROM[2168] <= 12'he89; 
SIN_ROM[2169] <= 12'he86; 
SIN_ROM[2170] <= 12'he83; 
SIN_ROM[2171] <= 12'he80; 
SIN_ROM[2172] <= 12'he7d; 
SIN_ROM[2173] <= 12'he7a; 
SIN_ROM[2174] <= 12'he77; 
SIN_ROM[2175] <= 12'he74; 
SIN_ROM[2176] <= 12'he71; 
SIN_ROM[2177] <= 12'he6e; 
SIN_ROM[2178] <= 12'he6a; 
SIN_ROM[2179] <= 12'he67; 
SIN_ROM[2180] <= 12'he64; 
SIN_ROM[2181] <= 12'he61; 
SIN_ROM[2182] <= 12'he5e; 
SIN_ROM[2183] <= 12'he5b; 
SIN_ROM[2184] <= 12'he58; 
SIN_ROM[2185] <= 12'he55; 
SIN_ROM[2186] <= 12'he52; 
SIN_ROM[2187] <= 12'he4f; 
SIN_ROM[2188] <= 12'he4c; 
SIN_ROM[2189] <= 12'he49; 
SIN_ROM[2190] <= 12'he46; 
SIN_ROM[2191] <= 12'he43; 
SIN_ROM[2192] <= 12'he3f; 
SIN_ROM[2193] <= 12'he3c; 
SIN_ROM[2194] <= 12'he39; 
SIN_ROM[2195] <= 12'he36; 
SIN_ROM[2196] <= 12'he33; 
SIN_ROM[2197] <= 12'he30; 
SIN_ROM[2198] <= 12'he2d; 
SIN_ROM[2199] <= 12'he2a; 
SIN_ROM[2200] <= 12'he27; 
SIN_ROM[2201] <= 12'he24; 
SIN_ROM[2202] <= 12'he21; 
SIN_ROM[2203] <= 12'he1e; 
SIN_ROM[2204] <= 12'he1b; 
SIN_ROM[2205] <= 12'he18; 
SIN_ROM[2206] <= 12'he15; 
SIN_ROM[2207] <= 12'he12; 
SIN_ROM[2208] <= 12'he0f; 
SIN_ROM[2209] <= 12'he0c; 
SIN_ROM[2210] <= 12'he09; 
SIN_ROM[2211] <= 12'he05; 
SIN_ROM[2212] <= 12'he02; 
SIN_ROM[2213] <= 12'hdff; 
SIN_ROM[2214] <= 12'hdfc; 
SIN_ROM[2215] <= 12'hdf9; 
SIN_ROM[2216] <= 12'hdf6; 
SIN_ROM[2217] <= 12'hdf3; 
SIN_ROM[2218] <= 12'hdf0; 
SIN_ROM[2219] <= 12'hded; 
SIN_ROM[2220] <= 12'hdea; 
SIN_ROM[2221] <= 12'hde7; 
SIN_ROM[2222] <= 12'hde4; 
SIN_ROM[2223] <= 12'hde1; 
SIN_ROM[2224] <= 12'hdde; 
SIN_ROM[2225] <= 12'hddb; 
SIN_ROM[2226] <= 12'hdd8; 
SIN_ROM[2227] <= 12'hdd5; 
SIN_ROM[2228] <= 12'hdd2; 
SIN_ROM[2229] <= 12'hdcf; 
SIN_ROM[2230] <= 12'hdcc; 
SIN_ROM[2231] <= 12'hdc9; 
SIN_ROM[2232] <= 12'hdc6; 
SIN_ROM[2233] <= 12'hdc3; 
SIN_ROM[2234] <= 12'hdc0; 
SIN_ROM[2235] <= 12'hdbd; 
SIN_ROM[2236] <= 12'hdba; 
SIN_ROM[2237] <= 12'hdb7; 
SIN_ROM[2238] <= 12'hdb4; 
SIN_ROM[2239] <= 12'hdb1; 
SIN_ROM[2240] <= 12'hdae; 
SIN_ROM[2241] <= 12'hdab; 
SIN_ROM[2242] <= 12'hda8; 
SIN_ROM[2243] <= 12'hda5; 
SIN_ROM[2244] <= 12'hda2; 
SIN_ROM[2245] <= 12'hd9f; 
SIN_ROM[2246] <= 12'hd9c; 
SIN_ROM[2247] <= 12'hd99; 
SIN_ROM[2248] <= 12'hd96; 
SIN_ROM[2249] <= 12'hd93; 
SIN_ROM[2250] <= 12'hd90; 
SIN_ROM[2251] <= 12'hd8d; 
SIN_ROM[2252] <= 12'hd8a; 
SIN_ROM[2253] <= 12'hd87; 
SIN_ROM[2254] <= 12'hd84; 
SIN_ROM[2255] <= 12'hd81; 
SIN_ROM[2256] <= 12'hd7e; 
SIN_ROM[2257] <= 12'hd7b; 
SIN_ROM[2258] <= 12'hd78; 
SIN_ROM[2259] <= 12'hd75; 
SIN_ROM[2260] <= 12'hd72; 
SIN_ROM[2261] <= 12'hd6f; 
SIN_ROM[2262] <= 12'hd6c; 
SIN_ROM[2263] <= 12'hd69; 
SIN_ROM[2264] <= 12'hd66; 
SIN_ROM[2265] <= 12'hd63; 
SIN_ROM[2266] <= 12'hd60; 
SIN_ROM[2267] <= 12'hd5d; 
SIN_ROM[2268] <= 12'hd5a; 
SIN_ROM[2269] <= 12'hd57; 
SIN_ROM[2270] <= 12'hd54; 
SIN_ROM[2271] <= 12'hd51; 
SIN_ROM[2272] <= 12'hd4e; 
SIN_ROM[2273] <= 12'hd4b; 
SIN_ROM[2274] <= 12'hd48; 
SIN_ROM[2275] <= 12'hd46; 
SIN_ROM[2276] <= 12'hd43; 
SIN_ROM[2277] <= 12'hd40; 
SIN_ROM[2278] <= 12'hd3d; 
SIN_ROM[2279] <= 12'hd3a; 
SIN_ROM[2280] <= 12'hd37; 
SIN_ROM[2281] <= 12'hd34; 
SIN_ROM[2282] <= 12'hd31; 
SIN_ROM[2283] <= 12'hd2e; 
SIN_ROM[2284] <= 12'hd2b; 
SIN_ROM[2285] <= 12'hd28; 
SIN_ROM[2286] <= 12'hd25; 
SIN_ROM[2287] <= 12'hd22; 
SIN_ROM[2288] <= 12'hd1f; 
SIN_ROM[2289] <= 12'hd1c; 
SIN_ROM[2290] <= 12'hd19; 
SIN_ROM[2291] <= 12'hd17; 
SIN_ROM[2292] <= 12'hd14; 
SIN_ROM[2293] <= 12'hd11; 
SIN_ROM[2294] <= 12'hd0e; 
SIN_ROM[2295] <= 12'hd0b; 
SIN_ROM[2296] <= 12'hd08; 
SIN_ROM[2297] <= 12'hd05; 
SIN_ROM[2298] <= 12'hd02; 
SIN_ROM[2299] <= 12'hcff; 
SIN_ROM[2300] <= 12'hcfc; 
SIN_ROM[2301] <= 12'hcf9; 
SIN_ROM[2302] <= 12'hcf6; 
SIN_ROM[2303] <= 12'hcf4; 
SIN_ROM[2304] <= 12'hcf1; 
SIN_ROM[2305] <= 12'hcee; 
SIN_ROM[2306] <= 12'hceb; 
SIN_ROM[2307] <= 12'hce8; 
SIN_ROM[2308] <= 12'hce5; 
SIN_ROM[2309] <= 12'hce2; 
SIN_ROM[2310] <= 12'hcdf; 
SIN_ROM[2311] <= 12'hcdc; 
SIN_ROM[2312] <= 12'hcd9; 
SIN_ROM[2313] <= 12'hcd7; 
SIN_ROM[2314] <= 12'hcd4; 
SIN_ROM[2315] <= 12'hcd1; 
SIN_ROM[2316] <= 12'hcce; 
SIN_ROM[2317] <= 12'hccb; 
SIN_ROM[2318] <= 12'hcc8; 
SIN_ROM[2319] <= 12'hcc5; 
SIN_ROM[2320] <= 12'hcc2; 
SIN_ROM[2321] <= 12'hcc0; 
SIN_ROM[2322] <= 12'hcbd; 
SIN_ROM[2323] <= 12'hcba; 
SIN_ROM[2324] <= 12'hcb7; 
SIN_ROM[2325] <= 12'hcb4; 
SIN_ROM[2326] <= 12'hcb1; 
SIN_ROM[2327] <= 12'hcae; 
SIN_ROM[2328] <= 12'hcac; 
SIN_ROM[2329] <= 12'hca9; 
SIN_ROM[2330] <= 12'hca6; 
SIN_ROM[2331] <= 12'hca3; 
SIN_ROM[2332] <= 12'hca0; 
SIN_ROM[2333] <= 12'hc9d; 
SIN_ROM[2334] <= 12'hc9a; 
SIN_ROM[2335] <= 12'hc98; 
SIN_ROM[2336] <= 12'hc95; 
SIN_ROM[2337] <= 12'hc92; 
SIN_ROM[2338] <= 12'hc8f; 
SIN_ROM[2339] <= 12'hc8c; 
SIN_ROM[2340] <= 12'hc89; 
SIN_ROM[2341] <= 12'hc87; 
SIN_ROM[2342] <= 12'hc84; 
SIN_ROM[2343] <= 12'hc81; 
SIN_ROM[2344] <= 12'hc7e; 
SIN_ROM[2345] <= 12'hc7b; 
SIN_ROM[2346] <= 12'hc79; 
SIN_ROM[2347] <= 12'hc76; 
SIN_ROM[2348] <= 12'hc73; 
SIN_ROM[2349] <= 12'hc70; 
SIN_ROM[2350] <= 12'hc6d; 
SIN_ROM[2351] <= 12'hc6a; 
SIN_ROM[2352] <= 12'hc68; 
SIN_ROM[2353] <= 12'hc65; 
SIN_ROM[2354] <= 12'hc62; 
SIN_ROM[2355] <= 12'hc5f; 
SIN_ROM[2356] <= 12'hc5c; 
SIN_ROM[2357] <= 12'hc5a; 
SIN_ROM[2358] <= 12'hc57; 
SIN_ROM[2359] <= 12'hc54; 
SIN_ROM[2360] <= 12'hc51; 
SIN_ROM[2361] <= 12'hc4e; 
SIN_ROM[2362] <= 12'hc4c; 
SIN_ROM[2363] <= 12'hc49; 
SIN_ROM[2364] <= 12'hc46; 
SIN_ROM[2365] <= 12'hc43; 
SIN_ROM[2366] <= 12'hc41; 
SIN_ROM[2367] <= 12'hc3e; 
SIN_ROM[2368] <= 12'hc3b; 
SIN_ROM[2369] <= 12'hc38; 
SIN_ROM[2370] <= 12'hc36; 
SIN_ROM[2371] <= 12'hc33; 
SIN_ROM[2372] <= 12'hc30; 
SIN_ROM[2373] <= 12'hc2d; 
SIN_ROM[2374] <= 12'hc2a; 
SIN_ROM[2375] <= 12'hc28; 
SIN_ROM[2376] <= 12'hc25; 
SIN_ROM[2377] <= 12'hc22; 
SIN_ROM[2378] <= 12'hc1f; 
SIN_ROM[2379] <= 12'hc1d; 
SIN_ROM[2380] <= 12'hc1a; 
SIN_ROM[2381] <= 12'hc17; 
SIN_ROM[2382] <= 12'hc15; 
SIN_ROM[2383] <= 12'hc12; 
SIN_ROM[2384] <= 12'hc0f; 
SIN_ROM[2385] <= 12'hc0c; 
SIN_ROM[2386] <= 12'hc0a; 
SIN_ROM[2387] <= 12'hc07; 
SIN_ROM[2388] <= 12'hc04; 
SIN_ROM[2389] <= 12'hc01; 
SIN_ROM[2390] <= 12'hbff; 
SIN_ROM[2391] <= 12'hbfc; 
SIN_ROM[2392] <= 12'hbf9; 
SIN_ROM[2393] <= 12'hbf7; 
SIN_ROM[2394] <= 12'hbf4; 
SIN_ROM[2395] <= 12'hbf1; 
SIN_ROM[2396] <= 12'hbee; 
SIN_ROM[2397] <= 12'hbec; 
SIN_ROM[2398] <= 12'hbe9; 
SIN_ROM[2399] <= 12'hbe6; 
SIN_ROM[2400] <= 12'hbe4; 
SIN_ROM[2401] <= 12'hbe1; 
SIN_ROM[2402] <= 12'hbde; 
SIN_ROM[2403] <= 12'hbdc; 
SIN_ROM[2404] <= 12'hbd9; 
SIN_ROM[2405] <= 12'hbd6; 
SIN_ROM[2406] <= 12'hbd4; 
SIN_ROM[2407] <= 12'hbd1; 
SIN_ROM[2408] <= 12'hbce; 
SIN_ROM[2409] <= 12'hbcb; 
SIN_ROM[2410] <= 12'hbc9; 
SIN_ROM[2411] <= 12'hbc6; 
SIN_ROM[2412] <= 12'hbc3; 
SIN_ROM[2413] <= 12'hbc1; 
SIN_ROM[2414] <= 12'hbbe; 
SIN_ROM[2415] <= 12'hbbc; 
SIN_ROM[2416] <= 12'hbb9; 
SIN_ROM[2417] <= 12'hbb6; 
SIN_ROM[2418] <= 12'hbb4; 
SIN_ROM[2419] <= 12'hbb1; 
SIN_ROM[2420] <= 12'hbae; 
SIN_ROM[2421] <= 12'hbac; 
SIN_ROM[2422] <= 12'hba9; 
SIN_ROM[2423] <= 12'hba6; 
SIN_ROM[2424] <= 12'hba4; 
SIN_ROM[2425] <= 12'hba1; 
SIN_ROM[2426] <= 12'hb9e; 
SIN_ROM[2427] <= 12'hb9c; 
SIN_ROM[2428] <= 12'hb99; 
SIN_ROM[2429] <= 12'hb97; 
SIN_ROM[2430] <= 12'hb94; 
SIN_ROM[2431] <= 12'hb91; 
SIN_ROM[2432] <= 12'hb8f; 
SIN_ROM[2433] <= 12'hb8c; 
SIN_ROM[2434] <= 12'hb8a; 
SIN_ROM[2435] <= 12'hb87; 
SIN_ROM[2436] <= 12'hb84; 
SIN_ROM[2437] <= 12'hb82; 
SIN_ROM[2438] <= 12'hb7f; 
SIN_ROM[2439] <= 12'hb7d; 
SIN_ROM[2440] <= 12'hb7a; 
SIN_ROM[2441] <= 12'hb77; 
SIN_ROM[2442] <= 12'hb75; 
SIN_ROM[2443] <= 12'hb72; 
SIN_ROM[2444] <= 12'hb70; 
SIN_ROM[2445] <= 12'hb6d; 
SIN_ROM[2446] <= 12'hb6a; 
SIN_ROM[2447] <= 12'hb68; 
SIN_ROM[2448] <= 12'hb65; 
SIN_ROM[2449] <= 12'hb63; 
SIN_ROM[2450] <= 12'hb60; 
SIN_ROM[2451] <= 12'hb5e; 
SIN_ROM[2452] <= 12'hb5b; 
SIN_ROM[2453] <= 12'hb59; 
SIN_ROM[2454] <= 12'hb56; 
SIN_ROM[2455] <= 12'hb53; 
SIN_ROM[2456] <= 12'hb51; 
SIN_ROM[2457] <= 12'hb4e; 
SIN_ROM[2458] <= 12'hb4c; 
SIN_ROM[2459] <= 12'hb49; 
SIN_ROM[2460] <= 12'hb47; 
SIN_ROM[2461] <= 12'hb44; 
SIN_ROM[2462] <= 12'hb42; 
SIN_ROM[2463] <= 12'hb3f; 
SIN_ROM[2464] <= 12'hb3d; 
SIN_ROM[2465] <= 12'hb3a; 
SIN_ROM[2466] <= 12'hb38; 
SIN_ROM[2467] <= 12'hb35; 
SIN_ROM[2468] <= 12'hb33; 
SIN_ROM[2469] <= 12'hb30; 
SIN_ROM[2470] <= 12'hb2e; 
SIN_ROM[2471] <= 12'hb2b; 
SIN_ROM[2472] <= 12'hb29; 
SIN_ROM[2473] <= 12'hb26; 
SIN_ROM[2474] <= 12'hb24; 
SIN_ROM[2475] <= 12'hb21; 
SIN_ROM[2476] <= 12'hb1f; 
SIN_ROM[2477] <= 12'hb1c; 
SIN_ROM[2478] <= 12'hb1a; 
SIN_ROM[2479] <= 12'hb17; 
SIN_ROM[2480] <= 12'hb15; 
SIN_ROM[2481] <= 12'hb12; 
SIN_ROM[2482] <= 12'hb10; 
SIN_ROM[2483] <= 12'hb0d; 
SIN_ROM[2484] <= 12'hb0b; 
SIN_ROM[2485] <= 12'hb08; 
SIN_ROM[2486] <= 12'hb06; 
SIN_ROM[2487] <= 12'hb03; 
SIN_ROM[2488] <= 12'hb01; 
SIN_ROM[2489] <= 12'hafe; 
SIN_ROM[2490] <= 12'hafc; 
SIN_ROM[2491] <= 12'hafa; 
SIN_ROM[2492] <= 12'haf7; 
SIN_ROM[2493] <= 12'haf5; 
SIN_ROM[2494] <= 12'haf2; 
SIN_ROM[2495] <= 12'haf0; 
SIN_ROM[2496] <= 12'haed; 
SIN_ROM[2497] <= 12'haeb; 
SIN_ROM[2498] <= 12'hae9; 
SIN_ROM[2499] <= 12'hae6; 
SIN_ROM[2500] <= 12'hae4; 
SIN_ROM[2501] <= 12'hae1; 
SIN_ROM[2502] <= 12'hadf; 
SIN_ROM[2503] <= 12'hadc; 
SIN_ROM[2504] <= 12'hada; 
SIN_ROM[2505] <= 12'had8; 
SIN_ROM[2506] <= 12'had5; 
SIN_ROM[2507] <= 12'had3; 
SIN_ROM[2508] <= 12'had0; 
SIN_ROM[2509] <= 12'hace; 
SIN_ROM[2510] <= 12'hacc; 
SIN_ROM[2511] <= 12'hac9; 
SIN_ROM[2512] <= 12'hac7; 
SIN_ROM[2513] <= 12'hac5; 
SIN_ROM[2514] <= 12'hac2; 
SIN_ROM[2515] <= 12'hac0; 
SIN_ROM[2516] <= 12'habd; 
SIN_ROM[2517] <= 12'habb; 
SIN_ROM[2518] <= 12'hab9; 
SIN_ROM[2519] <= 12'hab6; 
SIN_ROM[2520] <= 12'hab4; 
SIN_ROM[2521] <= 12'hab2; 
SIN_ROM[2522] <= 12'haaf; 
SIN_ROM[2523] <= 12'haad; 
SIN_ROM[2524] <= 12'haab; 
SIN_ROM[2525] <= 12'haa8; 
SIN_ROM[2526] <= 12'haa6; 
SIN_ROM[2527] <= 12'haa4; 
SIN_ROM[2528] <= 12'haa1; 
SIN_ROM[2529] <= 12'ha9f; 
SIN_ROM[2530] <= 12'ha9d; 
SIN_ROM[2531] <= 12'ha9a; 
SIN_ROM[2532] <= 12'ha98; 
SIN_ROM[2533] <= 12'ha96; 
SIN_ROM[2534] <= 12'ha93; 
SIN_ROM[2535] <= 12'ha91; 
SIN_ROM[2536] <= 12'ha8f; 
SIN_ROM[2537] <= 12'ha8d; 
SIN_ROM[2538] <= 12'ha8a; 
SIN_ROM[2539] <= 12'ha88; 
SIN_ROM[2540] <= 12'ha86; 
SIN_ROM[2541] <= 12'ha83; 
SIN_ROM[2542] <= 12'ha81; 
SIN_ROM[2543] <= 12'ha7f; 
SIN_ROM[2544] <= 12'ha7d; 
SIN_ROM[2545] <= 12'ha7a; 
SIN_ROM[2546] <= 12'ha78; 
SIN_ROM[2547] <= 12'ha76; 
SIN_ROM[2548] <= 12'ha73; 
SIN_ROM[2549] <= 12'ha71; 
SIN_ROM[2550] <= 12'ha6f; 
SIN_ROM[2551] <= 12'ha6d; 
SIN_ROM[2552] <= 12'ha6a; 
SIN_ROM[2553] <= 12'ha68; 
SIN_ROM[2554] <= 12'ha66; 
SIN_ROM[2555] <= 12'ha64; 
SIN_ROM[2556] <= 12'ha61; 
SIN_ROM[2557] <= 12'ha5f; 
SIN_ROM[2558] <= 12'ha5d; 
SIN_ROM[2559] <= 12'ha5b; 
SIN_ROM[2560] <= 12'ha59; 
SIN_ROM[2561] <= 12'ha56; 
SIN_ROM[2562] <= 12'ha54; 
SIN_ROM[2563] <= 12'ha52; 
SIN_ROM[2564] <= 12'ha50; 
SIN_ROM[2565] <= 12'ha4d; 
SIN_ROM[2566] <= 12'ha4b; 
SIN_ROM[2567] <= 12'ha49; 
SIN_ROM[2568] <= 12'ha47; 
SIN_ROM[2569] <= 12'ha45; 
SIN_ROM[2570] <= 12'ha43; 
SIN_ROM[2571] <= 12'ha40; 
SIN_ROM[2572] <= 12'ha3e; 
SIN_ROM[2573] <= 12'ha3c; 
SIN_ROM[2574] <= 12'ha3a; 
SIN_ROM[2575] <= 12'ha38; 
SIN_ROM[2576] <= 12'ha35; 
SIN_ROM[2577] <= 12'ha33; 
SIN_ROM[2578] <= 12'ha31; 
SIN_ROM[2579] <= 12'ha2f; 
SIN_ROM[2580] <= 12'ha2d; 
SIN_ROM[2581] <= 12'ha2b; 
SIN_ROM[2582] <= 12'ha29; 
SIN_ROM[2583] <= 12'ha26; 
SIN_ROM[2584] <= 12'ha24; 
SIN_ROM[2585] <= 12'ha22; 
SIN_ROM[2586] <= 12'ha20; 
SIN_ROM[2587] <= 12'ha1e; 
SIN_ROM[2588] <= 12'ha1c; 
SIN_ROM[2589] <= 12'ha1a; 
SIN_ROM[2590] <= 12'ha17; 
SIN_ROM[2591] <= 12'ha15; 
SIN_ROM[2592] <= 12'ha13; 
SIN_ROM[2593] <= 12'ha11; 
SIN_ROM[2594] <= 12'ha0f; 
SIN_ROM[2595] <= 12'ha0d; 
SIN_ROM[2596] <= 12'ha0b; 
SIN_ROM[2597] <= 12'ha09; 
SIN_ROM[2598] <= 12'ha07; 
SIN_ROM[2599] <= 12'ha05; 
SIN_ROM[2600] <= 12'ha03; 
SIN_ROM[2601] <= 12'ha00; 
SIN_ROM[2602] <= 12'h9fe; 
SIN_ROM[2603] <= 12'h9fc; 
SIN_ROM[2604] <= 12'h9fa; 
SIN_ROM[2605] <= 12'h9f8; 
SIN_ROM[2606] <= 12'h9f6; 
SIN_ROM[2607] <= 12'h9f4; 
SIN_ROM[2608] <= 12'h9f2; 
SIN_ROM[2609] <= 12'h9f0; 
SIN_ROM[2610] <= 12'h9ee; 
SIN_ROM[2611] <= 12'h9ec; 
SIN_ROM[2612] <= 12'h9ea; 
SIN_ROM[2613] <= 12'h9e8; 
SIN_ROM[2614] <= 12'h9e6; 
SIN_ROM[2615] <= 12'h9e4; 
SIN_ROM[2616] <= 12'h9e2; 
SIN_ROM[2617] <= 12'h9e0; 
SIN_ROM[2618] <= 12'h9de; 
SIN_ROM[2619] <= 12'h9dc; 
SIN_ROM[2620] <= 12'h9da; 
SIN_ROM[2621] <= 12'h9d8; 
SIN_ROM[2622] <= 12'h9d6; 
SIN_ROM[2623] <= 12'h9d4; 
SIN_ROM[2624] <= 12'h9d2; 
SIN_ROM[2625] <= 12'h9d0; 
SIN_ROM[2626] <= 12'h9ce; 
SIN_ROM[2627] <= 12'h9cc; 
SIN_ROM[2628] <= 12'h9ca; 
SIN_ROM[2629] <= 12'h9c8; 
SIN_ROM[2630] <= 12'h9c6; 
SIN_ROM[2631] <= 12'h9c4; 
SIN_ROM[2632] <= 12'h9c2; 
SIN_ROM[2633] <= 12'h9c0; 
SIN_ROM[2634] <= 12'h9be; 
SIN_ROM[2635] <= 12'h9bc; 
SIN_ROM[2636] <= 12'h9ba; 
SIN_ROM[2637] <= 12'h9b8; 
SIN_ROM[2638] <= 12'h9b6; 
SIN_ROM[2639] <= 12'h9b4; 
SIN_ROM[2640] <= 12'h9b2; 
SIN_ROM[2641] <= 12'h9b0; 
SIN_ROM[2642] <= 12'h9ae; 
SIN_ROM[2643] <= 12'h9ac; 
SIN_ROM[2644] <= 12'h9ab; 
SIN_ROM[2645] <= 12'h9a9; 
SIN_ROM[2646] <= 12'h9a7; 
SIN_ROM[2647] <= 12'h9a5; 
SIN_ROM[2648] <= 12'h9a3; 
SIN_ROM[2649] <= 12'h9a1; 
SIN_ROM[2650] <= 12'h99f; 
SIN_ROM[2651] <= 12'h99d; 
SIN_ROM[2652] <= 12'h99b; 
SIN_ROM[2653] <= 12'h999; 
SIN_ROM[2654] <= 12'h998; 
SIN_ROM[2655] <= 12'h996; 
SIN_ROM[2656] <= 12'h994; 
SIN_ROM[2657] <= 12'h992; 
SIN_ROM[2658] <= 12'h990; 
SIN_ROM[2659] <= 12'h98e; 
SIN_ROM[2660] <= 12'h98c; 
SIN_ROM[2661] <= 12'h98b; 
SIN_ROM[2662] <= 12'h989; 
SIN_ROM[2663] <= 12'h987; 
SIN_ROM[2664] <= 12'h985; 
SIN_ROM[2665] <= 12'h983; 
SIN_ROM[2666] <= 12'h981; 
SIN_ROM[2667] <= 12'h97f; 
SIN_ROM[2668] <= 12'h97e; 
SIN_ROM[2669] <= 12'h97c; 
SIN_ROM[2670] <= 12'h97a; 
SIN_ROM[2671] <= 12'h978; 
SIN_ROM[2672] <= 12'h976; 
SIN_ROM[2673] <= 12'h975; 
SIN_ROM[2674] <= 12'h973; 
SIN_ROM[2675] <= 12'h971; 
SIN_ROM[2676] <= 12'h96f; 
SIN_ROM[2677] <= 12'h96d; 
SIN_ROM[2678] <= 12'h96c; 
SIN_ROM[2679] <= 12'h96a; 
SIN_ROM[2680] <= 12'h968; 
SIN_ROM[2681] <= 12'h966; 
SIN_ROM[2682] <= 12'h965; 
SIN_ROM[2683] <= 12'h963; 
SIN_ROM[2684] <= 12'h961; 
SIN_ROM[2685] <= 12'h95f; 
SIN_ROM[2686] <= 12'h95d; 
SIN_ROM[2687] <= 12'h95c; 
SIN_ROM[2688] <= 12'h95a; 
SIN_ROM[2689] <= 12'h958; 
SIN_ROM[2690] <= 12'h957; 
SIN_ROM[2691] <= 12'h955; 
SIN_ROM[2692] <= 12'h953; 
SIN_ROM[2693] <= 12'h951; 
SIN_ROM[2694] <= 12'h950; 
SIN_ROM[2695] <= 12'h94e; 
SIN_ROM[2696] <= 12'h94c; 
SIN_ROM[2697] <= 12'h94a; 
SIN_ROM[2698] <= 12'h949; 
SIN_ROM[2699] <= 12'h947; 
SIN_ROM[2700] <= 12'h945; 
SIN_ROM[2701] <= 12'h944; 
SIN_ROM[2702] <= 12'h942; 
SIN_ROM[2703] <= 12'h940; 
SIN_ROM[2704] <= 12'h93f; 
SIN_ROM[2705] <= 12'h93d; 
SIN_ROM[2706] <= 12'h93b; 
SIN_ROM[2707] <= 12'h93a; 
SIN_ROM[2708] <= 12'h938; 
SIN_ROM[2709] <= 12'h936; 
SIN_ROM[2710] <= 12'h935; 
SIN_ROM[2711] <= 12'h933; 
SIN_ROM[2712] <= 12'h931; 
SIN_ROM[2713] <= 12'h930; 
SIN_ROM[2714] <= 12'h92e; 
SIN_ROM[2715] <= 12'h92c; 
SIN_ROM[2716] <= 12'h92b; 
SIN_ROM[2717] <= 12'h929; 
SIN_ROM[2718] <= 12'h927; 
SIN_ROM[2719] <= 12'h926; 
SIN_ROM[2720] <= 12'h924; 
SIN_ROM[2721] <= 12'h923; 
SIN_ROM[2722] <= 12'h921; 
SIN_ROM[2723] <= 12'h91f; 
SIN_ROM[2724] <= 12'h91e; 
SIN_ROM[2725] <= 12'h91c; 
SIN_ROM[2726] <= 12'h91b; 
SIN_ROM[2727] <= 12'h919; 
SIN_ROM[2728] <= 12'h917; 
SIN_ROM[2729] <= 12'h916; 
SIN_ROM[2730] <= 12'h914; 
SIN_ROM[2731] <= 12'h913; 
SIN_ROM[2732] <= 12'h911; 
SIN_ROM[2733] <= 12'h910; 
SIN_ROM[2734] <= 12'h90e; 
SIN_ROM[2735] <= 12'h90c; 
SIN_ROM[2736] <= 12'h90b; 
SIN_ROM[2737] <= 12'h909; 
SIN_ROM[2738] <= 12'h908; 
SIN_ROM[2739] <= 12'h906; 
SIN_ROM[2740] <= 12'h905; 
SIN_ROM[2741] <= 12'h903; 
SIN_ROM[2742] <= 12'h902; 
SIN_ROM[2743] <= 12'h900; 
SIN_ROM[2744] <= 12'h8ff; 
SIN_ROM[2745] <= 12'h8fd; 
SIN_ROM[2746] <= 12'h8fc; 
SIN_ROM[2747] <= 12'h8fa; 
SIN_ROM[2748] <= 12'h8f9; 
SIN_ROM[2749] <= 12'h8f7; 
SIN_ROM[2750] <= 12'h8f6; 
SIN_ROM[2751] <= 12'h8f4; 
SIN_ROM[2752] <= 12'h8f3; 
SIN_ROM[2753] <= 12'h8f1; 
SIN_ROM[2754] <= 12'h8f0; 
SIN_ROM[2755] <= 12'h8ee; 
SIN_ROM[2756] <= 12'h8ed; 
SIN_ROM[2757] <= 12'h8eb; 
SIN_ROM[2758] <= 12'h8ea; 
SIN_ROM[2759] <= 12'h8e8; 
SIN_ROM[2760] <= 12'h8e7; 
SIN_ROM[2761] <= 12'h8e6; 
SIN_ROM[2762] <= 12'h8e4; 
SIN_ROM[2763] <= 12'h8e3; 
SIN_ROM[2764] <= 12'h8e1; 
SIN_ROM[2765] <= 12'h8e0; 
SIN_ROM[2766] <= 12'h8de; 
SIN_ROM[2767] <= 12'h8dd; 
SIN_ROM[2768] <= 12'h8dc; 
SIN_ROM[2769] <= 12'h8da; 
SIN_ROM[2770] <= 12'h8d9; 
SIN_ROM[2771] <= 12'h8d7; 
SIN_ROM[2772] <= 12'h8d6; 
SIN_ROM[2773] <= 12'h8d5; 
SIN_ROM[2774] <= 12'h8d3; 
SIN_ROM[2775] <= 12'h8d2; 
SIN_ROM[2776] <= 12'h8d0; 
SIN_ROM[2777] <= 12'h8cf; 
SIN_ROM[2778] <= 12'h8ce; 
SIN_ROM[2779] <= 12'h8cc; 
SIN_ROM[2780] <= 12'h8cb; 
SIN_ROM[2781] <= 12'h8ca; 
SIN_ROM[2782] <= 12'h8c8; 
SIN_ROM[2783] <= 12'h8c7; 
SIN_ROM[2784] <= 12'h8c6; 
SIN_ROM[2785] <= 12'h8c4; 
SIN_ROM[2786] <= 12'h8c3; 
SIN_ROM[2787] <= 12'h8c2; 
SIN_ROM[2788] <= 12'h8c0; 
SIN_ROM[2789] <= 12'h8bf; 
SIN_ROM[2790] <= 12'h8be; 
SIN_ROM[2791] <= 12'h8bc; 
SIN_ROM[2792] <= 12'h8bb; 
SIN_ROM[2793] <= 12'h8ba; 
SIN_ROM[2794] <= 12'h8b8; 
SIN_ROM[2795] <= 12'h8b7; 
SIN_ROM[2796] <= 12'h8b6; 
SIN_ROM[2797] <= 12'h8b4; 
SIN_ROM[2798] <= 12'h8b3; 
SIN_ROM[2799] <= 12'h8b2; 
SIN_ROM[2800] <= 12'h8b1; 
SIN_ROM[2801] <= 12'h8af; 
SIN_ROM[2802] <= 12'h8ae; 
SIN_ROM[2803] <= 12'h8ad; 
SIN_ROM[2804] <= 12'h8ac; 
SIN_ROM[2805] <= 12'h8aa; 
SIN_ROM[2806] <= 12'h8a9; 
SIN_ROM[2807] <= 12'h8a8; 
SIN_ROM[2808] <= 12'h8a7; 
SIN_ROM[2809] <= 12'h8a5; 
SIN_ROM[2810] <= 12'h8a4; 
SIN_ROM[2811] <= 12'h8a3; 
SIN_ROM[2812] <= 12'h8a2; 
SIN_ROM[2813] <= 12'h8a0; 
SIN_ROM[2814] <= 12'h89f; 
SIN_ROM[2815] <= 12'h89e; 
SIN_ROM[2816] <= 12'h89d; 
SIN_ROM[2817] <= 12'h89c; 
SIN_ROM[2818] <= 12'h89a; 
SIN_ROM[2819] <= 12'h899; 
SIN_ROM[2820] <= 12'h898; 
SIN_ROM[2821] <= 12'h897; 
SIN_ROM[2822] <= 12'h896; 
SIN_ROM[2823] <= 12'h895; 
SIN_ROM[2824] <= 12'h893; 
SIN_ROM[2825] <= 12'h892; 
SIN_ROM[2826] <= 12'h891; 
SIN_ROM[2827] <= 12'h890; 
SIN_ROM[2828] <= 12'h88f; 
SIN_ROM[2829] <= 12'h88e; 
SIN_ROM[2830] <= 12'h88c; 
SIN_ROM[2831] <= 12'h88b; 
SIN_ROM[2832] <= 12'h88a; 
SIN_ROM[2833] <= 12'h889; 
SIN_ROM[2834] <= 12'h888; 
SIN_ROM[2835] <= 12'h887; 
SIN_ROM[2836] <= 12'h886; 
SIN_ROM[2837] <= 12'h885; 
SIN_ROM[2838] <= 12'h883; 
SIN_ROM[2839] <= 12'h882; 
SIN_ROM[2840] <= 12'h881; 
SIN_ROM[2841] <= 12'h880; 
SIN_ROM[2842] <= 12'h87f; 
SIN_ROM[2843] <= 12'h87e; 
SIN_ROM[2844] <= 12'h87d; 
SIN_ROM[2845] <= 12'h87c; 
SIN_ROM[2846] <= 12'h87b; 
SIN_ROM[2847] <= 12'h87a; 
SIN_ROM[2848] <= 12'h879; 
SIN_ROM[2849] <= 12'h878; 
SIN_ROM[2850] <= 12'h877; 
SIN_ROM[2851] <= 12'h876; 
SIN_ROM[2852] <= 12'h874; 
SIN_ROM[2853] <= 12'h873; 
SIN_ROM[2854] <= 12'h872; 
SIN_ROM[2855] <= 12'h871; 
SIN_ROM[2856] <= 12'h870; 
SIN_ROM[2857] <= 12'h86f; 
SIN_ROM[2858] <= 12'h86e; 
SIN_ROM[2859] <= 12'h86d; 
SIN_ROM[2860] <= 12'h86c; 
SIN_ROM[2861] <= 12'h86b; 
SIN_ROM[2862] <= 12'h86a; 
SIN_ROM[2863] <= 12'h869; 
SIN_ROM[2864] <= 12'h868; 
SIN_ROM[2865] <= 12'h867; 
SIN_ROM[2866] <= 12'h866; 
SIN_ROM[2867] <= 12'h865; 
SIN_ROM[2868] <= 12'h864; 
SIN_ROM[2869] <= 12'h863; 
SIN_ROM[2870] <= 12'h862; 
SIN_ROM[2871] <= 12'h862; 
SIN_ROM[2872] <= 12'h861; 
SIN_ROM[2873] <= 12'h860; 
SIN_ROM[2874] <= 12'h85f; 
SIN_ROM[2875] <= 12'h85e; 
SIN_ROM[2876] <= 12'h85d; 
SIN_ROM[2877] <= 12'h85c; 
SIN_ROM[2878] <= 12'h85b; 
SIN_ROM[2879] <= 12'h85a; 
SIN_ROM[2880] <= 12'h859; 
SIN_ROM[2881] <= 12'h858; 
SIN_ROM[2882] <= 12'h857; 
SIN_ROM[2883] <= 12'h856; 
SIN_ROM[2884] <= 12'h856; 
SIN_ROM[2885] <= 12'h855; 
SIN_ROM[2886] <= 12'h854; 
SIN_ROM[2887] <= 12'h853; 
SIN_ROM[2888] <= 12'h852; 
SIN_ROM[2889] <= 12'h851; 
SIN_ROM[2890] <= 12'h850; 
SIN_ROM[2891] <= 12'h84f; 
SIN_ROM[2892] <= 12'h84f; 
SIN_ROM[2893] <= 12'h84e; 
SIN_ROM[2894] <= 12'h84d; 
SIN_ROM[2895] <= 12'h84c; 
SIN_ROM[2896] <= 12'h84b; 
SIN_ROM[2897] <= 12'h84a; 
SIN_ROM[2898] <= 12'h849; 
SIN_ROM[2899] <= 12'h849; 
SIN_ROM[2900] <= 12'h848; 
SIN_ROM[2901] <= 12'h847; 
SIN_ROM[2902] <= 12'h846; 
SIN_ROM[2903] <= 12'h845; 
SIN_ROM[2904] <= 12'h845; 
SIN_ROM[2905] <= 12'h844; 
SIN_ROM[2906] <= 12'h843; 
SIN_ROM[2907] <= 12'h842; 
SIN_ROM[2908] <= 12'h841; 
SIN_ROM[2909] <= 12'h841; 
SIN_ROM[2910] <= 12'h840; 
SIN_ROM[2911] <= 12'h83f; 
SIN_ROM[2912] <= 12'h83e; 
SIN_ROM[2913] <= 12'h83e; 
SIN_ROM[2914] <= 12'h83d; 
SIN_ROM[2915] <= 12'h83c; 
SIN_ROM[2916] <= 12'h83b; 
SIN_ROM[2917] <= 12'h83b; 
SIN_ROM[2918] <= 12'h83a; 
SIN_ROM[2919] <= 12'h839; 
SIN_ROM[2920] <= 12'h838; 
SIN_ROM[2921] <= 12'h838; 
SIN_ROM[2922] <= 12'h837; 
SIN_ROM[2923] <= 12'h836; 
SIN_ROM[2924] <= 12'h836; 
SIN_ROM[2925] <= 12'h835; 
SIN_ROM[2926] <= 12'h834; 
SIN_ROM[2927] <= 12'h833; 
SIN_ROM[2928] <= 12'h833; 
SIN_ROM[2929] <= 12'h832; 
SIN_ROM[2930] <= 12'h831; 
SIN_ROM[2931] <= 12'h831; 
SIN_ROM[2932] <= 12'h830; 
SIN_ROM[2933] <= 12'h82f; 
SIN_ROM[2934] <= 12'h82f; 
SIN_ROM[2935] <= 12'h82e; 
SIN_ROM[2936] <= 12'h82d; 
SIN_ROM[2937] <= 12'h82d; 
SIN_ROM[2938] <= 12'h82c; 
SIN_ROM[2939] <= 12'h82b; 
SIN_ROM[2940] <= 12'h82b; 
SIN_ROM[2941] <= 12'h82a; 
SIN_ROM[2942] <= 12'h82a; 
SIN_ROM[2943] <= 12'h829; 
SIN_ROM[2944] <= 12'h828; 
SIN_ROM[2945] <= 12'h828; 
SIN_ROM[2946] <= 12'h827; 
SIN_ROM[2947] <= 12'h827; 
SIN_ROM[2948] <= 12'h826; 
SIN_ROM[2949] <= 12'h825; 
SIN_ROM[2950] <= 12'h825; 
SIN_ROM[2951] <= 12'h824; 
SIN_ROM[2952] <= 12'h824; 
SIN_ROM[2953] <= 12'h823; 
SIN_ROM[2954] <= 12'h822; 
SIN_ROM[2955] <= 12'h822; 
SIN_ROM[2956] <= 12'h821; 
SIN_ROM[2957] <= 12'h821; 
SIN_ROM[2958] <= 12'h820; 
SIN_ROM[2959] <= 12'h820; 
SIN_ROM[2960] <= 12'h81f; 
SIN_ROM[2961] <= 12'h81f; 
SIN_ROM[2962] <= 12'h81e; 
SIN_ROM[2963] <= 12'h81e; 
SIN_ROM[2964] <= 12'h81d; 
SIN_ROM[2965] <= 12'h81d; 
SIN_ROM[2966] <= 12'h81c; 
SIN_ROM[2967] <= 12'h81b; 
SIN_ROM[2968] <= 12'h81b; 
SIN_ROM[2969] <= 12'h81a; 
SIN_ROM[2970] <= 12'h81a; 
SIN_ROM[2971] <= 12'h81a; 
SIN_ROM[2972] <= 12'h819; 
SIN_ROM[2973] <= 12'h819; 
SIN_ROM[2974] <= 12'h818; 
SIN_ROM[2975] <= 12'h818; 
SIN_ROM[2976] <= 12'h817; 
SIN_ROM[2977] <= 12'h817; 
SIN_ROM[2978] <= 12'h816; 
SIN_ROM[2979] <= 12'h816; 
SIN_ROM[2980] <= 12'h815; 
SIN_ROM[2981] <= 12'h815; 
SIN_ROM[2982] <= 12'h814; 
SIN_ROM[2983] <= 12'h814; 
SIN_ROM[2984] <= 12'h814; 
SIN_ROM[2985] <= 12'h813; 
SIN_ROM[2986] <= 12'h813; 
SIN_ROM[2987] <= 12'h812; 
SIN_ROM[2988] <= 12'h812; 
SIN_ROM[2989] <= 12'h812; 
SIN_ROM[2990] <= 12'h811; 
SIN_ROM[2991] <= 12'h811; 
SIN_ROM[2992] <= 12'h810; 
SIN_ROM[2993] <= 12'h810; 
SIN_ROM[2994] <= 12'h810; 
SIN_ROM[2995] <= 12'h80f; 
SIN_ROM[2996] <= 12'h80f; 
SIN_ROM[2997] <= 12'h80f; 
SIN_ROM[2998] <= 12'h80e; 
SIN_ROM[2999] <= 12'h80e; 
SIN_ROM[3000] <= 12'h80d; 
SIN_ROM[3001] <= 12'h80d; 
SIN_ROM[3002] <= 12'h80d; 
SIN_ROM[3003] <= 12'h80c; 
SIN_ROM[3004] <= 12'h80c; 
SIN_ROM[3005] <= 12'h80c; 
SIN_ROM[3006] <= 12'h80b; 
SIN_ROM[3007] <= 12'h80b; 
SIN_ROM[3008] <= 12'h80b; 
SIN_ROM[3009] <= 12'h80b; 
SIN_ROM[3010] <= 12'h80a; 
SIN_ROM[3011] <= 12'h80a; 
SIN_ROM[3012] <= 12'h80a; 
SIN_ROM[3013] <= 12'h809; 
SIN_ROM[3014] <= 12'h809; 
SIN_ROM[3015] <= 12'h809; 
SIN_ROM[3016] <= 12'h809; 
SIN_ROM[3017] <= 12'h808; 
SIN_ROM[3018] <= 12'h808; 
SIN_ROM[3019] <= 12'h808; 
SIN_ROM[3020] <= 12'h808; 
SIN_ROM[3021] <= 12'h807; 
SIN_ROM[3022] <= 12'h807; 
SIN_ROM[3023] <= 12'h807; 
SIN_ROM[3024] <= 12'h807; 
SIN_ROM[3025] <= 12'h806; 
SIN_ROM[3026] <= 12'h806; 
SIN_ROM[3027] <= 12'h806; 
SIN_ROM[3028] <= 12'h806; 
SIN_ROM[3029] <= 12'h805; 
SIN_ROM[3030] <= 12'h805; 
SIN_ROM[3031] <= 12'h805; 
SIN_ROM[3032] <= 12'h805; 
SIN_ROM[3033] <= 12'h805; 
SIN_ROM[3034] <= 12'h804; 
SIN_ROM[3035] <= 12'h804; 
SIN_ROM[3036] <= 12'h804; 
SIN_ROM[3037] <= 12'h804; 
SIN_ROM[3038] <= 12'h804; 
SIN_ROM[3039] <= 12'h804; 
SIN_ROM[3040] <= 12'h803; 
SIN_ROM[3041] <= 12'h803; 
SIN_ROM[3042] <= 12'h803; 
SIN_ROM[3043] <= 12'h803; 
SIN_ROM[3044] <= 12'h803; 
SIN_ROM[3045] <= 12'h803; 
SIN_ROM[3046] <= 12'h803; 
SIN_ROM[3047] <= 12'h803; 
SIN_ROM[3048] <= 12'h802; 
SIN_ROM[3049] <= 12'h802; 
SIN_ROM[3050] <= 12'h802; 
SIN_ROM[3051] <= 12'h802; 
SIN_ROM[3052] <= 12'h802; 
SIN_ROM[3053] <= 12'h802; 
SIN_ROM[3054] <= 12'h802; 
SIN_ROM[3055] <= 12'h802; 
SIN_ROM[3056] <= 12'h802; 
SIN_ROM[3057] <= 12'h802; 
SIN_ROM[3058] <= 12'h801; 
SIN_ROM[3059] <= 12'h801; 
SIN_ROM[3060] <= 12'h801; 
SIN_ROM[3061] <= 12'h801; 
SIN_ROM[3062] <= 12'h801; 
SIN_ROM[3063] <= 12'h801; 
SIN_ROM[3064] <= 12'h801; 
SIN_ROM[3065] <= 12'h801; 
SIN_ROM[3066] <= 12'h801; 
SIN_ROM[3067] <= 12'h801; 
SIN_ROM[3068] <= 12'h801; 
SIN_ROM[3069] <= 12'h801; 
SIN_ROM[3070] <= 12'h801; 
SIN_ROM[3071] <= 12'h801; 
SIN_ROM[3072] <= 12'h801; 
SIN_ROM[3073] <= 12'h801; 
SIN_ROM[3074] <= 12'h801; 
SIN_ROM[3075] <= 12'h801; 
SIN_ROM[3076] <= 12'h801; 
SIN_ROM[3077] <= 12'h801; 
SIN_ROM[3078] <= 12'h801; 
SIN_ROM[3079] <= 12'h801; 
SIN_ROM[3080] <= 12'h801; 
SIN_ROM[3081] <= 12'h801; 
SIN_ROM[3082] <= 12'h801; 
SIN_ROM[3083] <= 12'h801; 
SIN_ROM[3084] <= 12'h801; 
SIN_ROM[3085] <= 12'h801; 
SIN_ROM[3086] <= 12'h801; 
SIN_ROM[3087] <= 12'h802; 
SIN_ROM[3088] <= 12'h802; 
SIN_ROM[3089] <= 12'h802; 
SIN_ROM[3090] <= 12'h802; 
SIN_ROM[3091] <= 12'h802; 
SIN_ROM[3092] <= 12'h802; 
SIN_ROM[3093] <= 12'h802; 
SIN_ROM[3094] <= 12'h802; 
SIN_ROM[3095] <= 12'h802; 
SIN_ROM[3096] <= 12'h802; 
SIN_ROM[3097] <= 12'h803; 
SIN_ROM[3098] <= 12'h803; 
SIN_ROM[3099] <= 12'h803; 
SIN_ROM[3100] <= 12'h803; 
SIN_ROM[3101] <= 12'h803; 
SIN_ROM[3102] <= 12'h803; 
SIN_ROM[3103] <= 12'h803; 
SIN_ROM[3104] <= 12'h803; 
SIN_ROM[3105] <= 12'h804; 
SIN_ROM[3106] <= 12'h804; 
SIN_ROM[3107] <= 12'h804; 
SIN_ROM[3108] <= 12'h804; 
SIN_ROM[3109] <= 12'h804; 
SIN_ROM[3110] <= 12'h804; 
SIN_ROM[3111] <= 12'h805; 
SIN_ROM[3112] <= 12'h805; 
SIN_ROM[3113] <= 12'h805; 
SIN_ROM[3114] <= 12'h805; 
SIN_ROM[3115] <= 12'h805; 
SIN_ROM[3116] <= 12'h806; 
SIN_ROM[3117] <= 12'h806; 
SIN_ROM[3118] <= 12'h806; 
SIN_ROM[3119] <= 12'h806; 
SIN_ROM[3120] <= 12'h807; 
SIN_ROM[3121] <= 12'h807; 
SIN_ROM[3122] <= 12'h807; 
SIN_ROM[3123] <= 12'h807; 
SIN_ROM[3124] <= 12'h808; 
SIN_ROM[3125] <= 12'h808; 
SIN_ROM[3126] <= 12'h808; 
SIN_ROM[3127] <= 12'h808; 
SIN_ROM[3128] <= 12'h809; 
SIN_ROM[3129] <= 12'h809; 
SIN_ROM[3130] <= 12'h809; 
SIN_ROM[3131] <= 12'h809; 
SIN_ROM[3132] <= 12'h80a; 
SIN_ROM[3133] <= 12'h80a; 
SIN_ROM[3134] <= 12'h80a; 
SIN_ROM[3135] <= 12'h80b; 
SIN_ROM[3136] <= 12'h80b; 
SIN_ROM[3137] <= 12'h80b; 
SIN_ROM[3138] <= 12'h80b; 
SIN_ROM[3139] <= 12'h80c; 
SIN_ROM[3140] <= 12'h80c; 
SIN_ROM[3141] <= 12'h80c; 
SIN_ROM[3142] <= 12'h80d; 
SIN_ROM[3143] <= 12'h80d; 
SIN_ROM[3144] <= 12'h80d; 
SIN_ROM[3145] <= 12'h80e; 
SIN_ROM[3146] <= 12'h80e; 
SIN_ROM[3147] <= 12'h80f; 
SIN_ROM[3148] <= 12'h80f; 
SIN_ROM[3149] <= 12'h80f; 
SIN_ROM[3150] <= 12'h810; 
SIN_ROM[3151] <= 12'h810; 
SIN_ROM[3152] <= 12'h810; 
SIN_ROM[3153] <= 12'h811; 
SIN_ROM[3154] <= 12'h811; 
SIN_ROM[3155] <= 12'h812; 
SIN_ROM[3156] <= 12'h812; 
SIN_ROM[3157] <= 12'h812; 
SIN_ROM[3158] <= 12'h813; 
SIN_ROM[3159] <= 12'h813; 
SIN_ROM[3160] <= 12'h814; 
SIN_ROM[3161] <= 12'h814; 
SIN_ROM[3162] <= 12'h814; 
SIN_ROM[3163] <= 12'h815; 
SIN_ROM[3164] <= 12'h815; 
SIN_ROM[3165] <= 12'h816; 
SIN_ROM[3166] <= 12'h816; 
SIN_ROM[3167] <= 12'h817; 
SIN_ROM[3168] <= 12'h817; 
SIN_ROM[3169] <= 12'h818; 
SIN_ROM[3170] <= 12'h818; 
SIN_ROM[3171] <= 12'h819; 
SIN_ROM[3172] <= 12'h819; 
SIN_ROM[3173] <= 12'h81a; 
SIN_ROM[3174] <= 12'h81a; 
SIN_ROM[3175] <= 12'h81a; 
SIN_ROM[3176] <= 12'h81b; 
SIN_ROM[3177] <= 12'h81b; 
SIN_ROM[3178] <= 12'h81c; 
SIN_ROM[3179] <= 12'h81d; 
SIN_ROM[3180] <= 12'h81d; 
SIN_ROM[3181] <= 12'h81e; 
SIN_ROM[3182] <= 12'h81e; 
SIN_ROM[3183] <= 12'h81f; 
SIN_ROM[3184] <= 12'h81f; 
SIN_ROM[3185] <= 12'h820; 
SIN_ROM[3186] <= 12'h820; 
SIN_ROM[3187] <= 12'h821; 
SIN_ROM[3188] <= 12'h821; 
SIN_ROM[3189] <= 12'h822; 
SIN_ROM[3190] <= 12'h822; 
SIN_ROM[3191] <= 12'h823; 
SIN_ROM[3192] <= 12'h824; 
SIN_ROM[3193] <= 12'h824; 
SIN_ROM[3194] <= 12'h825; 
SIN_ROM[3195] <= 12'h825; 
SIN_ROM[3196] <= 12'h826; 
SIN_ROM[3197] <= 12'h827; 
SIN_ROM[3198] <= 12'h827; 
SIN_ROM[3199] <= 12'h828; 
SIN_ROM[3200] <= 12'h828; 
SIN_ROM[3201] <= 12'h829; 
SIN_ROM[3202] <= 12'h82a; 
SIN_ROM[3203] <= 12'h82a; 
SIN_ROM[3204] <= 12'h82b; 
SIN_ROM[3205] <= 12'h82b; 
SIN_ROM[3206] <= 12'h82c; 
SIN_ROM[3207] <= 12'h82d; 
SIN_ROM[3208] <= 12'h82d; 
SIN_ROM[3209] <= 12'h82e; 
SIN_ROM[3210] <= 12'h82f; 
SIN_ROM[3211] <= 12'h82f; 
SIN_ROM[3212] <= 12'h830; 
SIN_ROM[3213] <= 12'h831; 
SIN_ROM[3214] <= 12'h831; 
SIN_ROM[3215] <= 12'h832; 
SIN_ROM[3216] <= 12'h833; 
SIN_ROM[3217] <= 12'h833; 
SIN_ROM[3218] <= 12'h834; 
SIN_ROM[3219] <= 12'h835; 
SIN_ROM[3220] <= 12'h836; 
SIN_ROM[3221] <= 12'h836; 
SIN_ROM[3222] <= 12'h837; 
SIN_ROM[3223] <= 12'h838; 
SIN_ROM[3224] <= 12'h838; 
SIN_ROM[3225] <= 12'h839; 
SIN_ROM[3226] <= 12'h83a; 
SIN_ROM[3227] <= 12'h83b; 
SIN_ROM[3228] <= 12'h83b; 
SIN_ROM[3229] <= 12'h83c; 
SIN_ROM[3230] <= 12'h83d; 
SIN_ROM[3231] <= 12'h83e; 
SIN_ROM[3232] <= 12'h83e; 
SIN_ROM[3233] <= 12'h83f; 
SIN_ROM[3234] <= 12'h840; 
SIN_ROM[3235] <= 12'h841; 
SIN_ROM[3236] <= 12'h841; 
SIN_ROM[3237] <= 12'h842; 
SIN_ROM[3238] <= 12'h843; 
SIN_ROM[3239] <= 12'h844; 
SIN_ROM[3240] <= 12'h845; 
SIN_ROM[3241] <= 12'h845; 
SIN_ROM[3242] <= 12'h846; 
SIN_ROM[3243] <= 12'h847; 
SIN_ROM[3244] <= 12'h848; 
SIN_ROM[3245] <= 12'h849; 
SIN_ROM[3246] <= 12'h849; 
SIN_ROM[3247] <= 12'h84a; 
SIN_ROM[3248] <= 12'h84b; 
SIN_ROM[3249] <= 12'h84c; 
SIN_ROM[3250] <= 12'h84d; 
SIN_ROM[3251] <= 12'h84e; 
SIN_ROM[3252] <= 12'h84f; 
SIN_ROM[3253] <= 12'h84f; 
SIN_ROM[3254] <= 12'h850; 
SIN_ROM[3255] <= 12'h851; 
SIN_ROM[3256] <= 12'h852; 
SIN_ROM[3257] <= 12'h853; 
SIN_ROM[3258] <= 12'h854; 
SIN_ROM[3259] <= 12'h855; 
SIN_ROM[3260] <= 12'h856; 
SIN_ROM[3261] <= 12'h856; 
SIN_ROM[3262] <= 12'h857; 
SIN_ROM[3263] <= 12'h858; 
SIN_ROM[3264] <= 12'h859; 
SIN_ROM[3265] <= 12'h85a; 
SIN_ROM[3266] <= 12'h85b; 
SIN_ROM[3267] <= 12'h85c; 
SIN_ROM[3268] <= 12'h85d; 
SIN_ROM[3269] <= 12'h85e; 
SIN_ROM[3270] <= 12'h85f; 
SIN_ROM[3271] <= 12'h860; 
SIN_ROM[3272] <= 12'h861; 
SIN_ROM[3273] <= 12'h862; 
SIN_ROM[3274] <= 12'h862; 
SIN_ROM[3275] <= 12'h863; 
SIN_ROM[3276] <= 12'h864; 
SIN_ROM[3277] <= 12'h865; 
SIN_ROM[3278] <= 12'h866; 
SIN_ROM[3279] <= 12'h867; 
SIN_ROM[3280] <= 12'h868; 
SIN_ROM[3281] <= 12'h869; 
SIN_ROM[3282] <= 12'h86a; 
SIN_ROM[3283] <= 12'h86b; 
SIN_ROM[3284] <= 12'h86c; 
SIN_ROM[3285] <= 12'h86d; 
SIN_ROM[3286] <= 12'h86e; 
SIN_ROM[3287] <= 12'h86f; 
SIN_ROM[3288] <= 12'h870; 
SIN_ROM[3289] <= 12'h871; 
SIN_ROM[3290] <= 12'h872; 
SIN_ROM[3291] <= 12'h873; 
SIN_ROM[3292] <= 12'h874; 
SIN_ROM[3293] <= 12'h876; 
SIN_ROM[3294] <= 12'h877; 
SIN_ROM[3295] <= 12'h878; 
SIN_ROM[3296] <= 12'h879; 
SIN_ROM[3297] <= 12'h87a; 
SIN_ROM[3298] <= 12'h87b; 
SIN_ROM[3299] <= 12'h87c; 
SIN_ROM[3300] <= 12'h87d; 
SIN_ROM[3301] <= 12'h87e; 
SIN_ROM[3302] <= 12'h87f; 
SIN_ROM[3303] <= 12'h880; 
SIN_ROM[3304] <= 12'h881; 
SIN_ROM[3305] <= 12'h882; 
SIN_ROM[3306] <= 12'h883; 
SIN_ROM[3307] <= 12'h885; 
SIN_ROM[3308] <= 12'h886; 
SIN_ROM[3309] <= 12'h887; 
SIN_ROM[3310] <= 12'h888; 
SIN_ROM[3311] <= 12'h889; 
SIN_ROM[3312] <= 12'h88a; 
SIN_ROM[3313] <= 12'h88b; 
SIN_ROM[3314] <= 12'h88c; 
SIN_ROM[3315] <= 12'h88e; 
SIN_ROM[3316] <= 12'h88f; 
SIN_ROM[3317] <= 12'h890; 
SIN_ROM[3318] <= 12'h891; 
SIN_ROM[3319] <= 12'h892; 
SIN_ROM[3320] <= 12'h893; 
SIN_ROM[3321] <= 12'h895; 
SIN_ROM[3322] <= 12'h896; 
SIN_ROM[3323] <= 12'h897; 
SIN_ROM[3324] <= 12'h898; 
SIN_ROM[3325] <= 12'h899; 
SIN_ROM[3326] <= 12'h89a; 
SIN_ROM[3327] <= 12'h89c; 
SIN_ROM[3328] <= 12'h89d; 
SIN_ROM[3329] <= 12'h89e; 
SIN_ROM[3330] <= 12'h89f; 
SIN_ROM[3331] <= 12'h8a0; 
SIN_ROM[3332] <= 12'h8a2; 
SIN_ROM[3333] <= 12'h8a3; 
SIN_ROM[3334] <= 12'h8a4; 
SIN_ROM[3335] <= 12'h8a5; 
SIN_ROM[3336] <= 12'h8a7; 
SIN_ROM[3337] <= 12'h8a8; 
SIN_ROM[3338] <= 12'h8a9; 
SIN_ROM[3339] <= 12'h8aa; 
SIN_ROM[3340] <= 12'h8ac; 
SIN_ROM[3341] <= 12'h8ad; 
SIN_ROM[3342] <= 12'h8ae; 
SIN_ROM[3343] <= 12'h8af; 
SIN_ROM[3344] <= 12'h8b1; 
SIN_ROM[3345] <= 12'h8b2; 
SIN_ROM[3346] <= 12'h8b3; 
SIN_ROM[3347] <= 12'h8b4; 
SIN_ROM[3348] <= 12'h8b6; 
SIN_ROM[3349] <= 12'h8b7; 
SIN_ROM[3350] <= 12'h8b8; 
SIN_ROM[3351] <= 12'h8ba; 
SIN_ROM[3352] <= 12'h8bb; 
SIN_ROM[3353] <= 12'h8bc; 
SIN_ROM[3354] <= 12'h8be; 
SIN_ROM[3355] <= 12'h8bf; 
SIN_ROM[3356] <= 12'h8c0; 
SIN_ROM[3357] <= 12'h8c2; 
SIN_ROM[3358] <= 12'h8c3; 
SIN_ROM[3359] <= 12'h8c4; 
SIN_ROM[3360] <= 12'h8c6; 
SIN_ROM[3361] <= 12'h8c7; 
SIN_ROM[3362] <= 12'h8c8; 
SIN_ROM[3363] <= 12'h8ca; 
SIN_ROM[3364] <= 12'h8cb; 
SIN_ROM[3365] <= 12'h8cc; 
SIN_ROM[3366] <= 12'h8ce; 
SIN_ROM[3367] <= 12'h8cf; 
SIN_ROM[3368] <= 12'h8d0; 
SIN_ROM[3369] <= 12'h8d2; 
SIN_ROM[3370] <= 12'h8d3; 
SIN_ROM[3371] <= 12'h8d5; 
SIN_ROM[3372] <= 12'h8d6; 
SIN_ROM[3373] <= 12'h8d7; 
SIN_ROM[3374] <= 12'h8d9; 
SIN_ROM[3375] <= 12'h8da; 
SIN_ROM[3376] <= 12'h8dc; 
SIN_ROM[3377] <= 12'h8dd; 
SIN_ROM[3378] <= 12'h8de; 
SIN_ROM[3379] <= 12'h8e0; 
SIN_ROM[3380] <= 12'h8e1; 
SIN_ROM[3381] <= 12'h8e3; 
SIN_ROM[3382] <= 12'h8e4; 
SIN_ROM[3383] <= 12'h8e6; 
SIN_ROM[3384] <= 12'h8e7; 
SIN_ROM[3385] <= 12'h8e8; 
SIN_ROM[3386] <= 12'h8ea; 
SIN_ROM[3387] <= 12'h8eb; 
SIN_ROM[3388] <= 12'h8ed; 
SIN_ROM[3389] <= 12'h8ee; 
SIN_ROM[3390] <= 12'h8f0; 
SIN_ROM[3391] <= 12'h8f1; 
SIN_ROM[3392] <= 12'h8f3; 
SIN_ROM[3393] <= 12'h8f4; 
SIN_ROM[3394] <= 12'h8f6; 
SIN_ROM[3395] <= 12'h8f7; 
SIN_ROM[3396] <= 12'h8f9; 
SIN_ROM[3397] <= 12'h8fa; 
SIN_ROM[3398] <= 12'h8fc; 
SIN_ROM[3399] <= 12'h8fd; 
SIN_ROM[3400] <= 12'h8ff; 
SIN_ROM[3401] <= 12'h900; 
SIN_ROM[3402] <= 12'h902; 
SIN_ROM[3403] <= 12'h903; 
SIN_ROM[3404] <= 12'h905; 
SIN_ROM[3405] <= 12'h906; 
SIN_ROM[3406] <= 12'h908; 
SIN_ROM[3407] <= 12'h909; 
SIN_ROM[3408] <= 12'h90b; 
SIN_ROM[3409] <= 12'h90c; 
SIN_ROM[3410] <= 12'h90e; 
SIN_ROM[3411] <= 12'h910; 
SIN_ROM[3412] <= 12'h911; 
SIN_ROM[3413] <= 12'h913; 
SIN_ROM[3414] <= 12'h914; 
SIN_ROM[3415] <= 12'h916; 
SIN_ROM[3416] <= 12'h917; 
SIN_ROM[3417] <= 12'h919; 
SIN_ROM[3418] <= 12'h91b; 
SIN_ROM[3419] <= 12'h91c; 
SIN_ROM[3420] <= 12'h91e; 
SIN_ROM[3421] <= 12'h91f; 
SIN_ROM[3422] <= 12'h921; 
SIN_ROM[3423] <= 12'h923; 
SIN_ROM[3424] <= 12'h924; 
SIN_ROM[3425] <= 12'h926; 
SIN_ROM[3426] <= 12'h927; 
SIN_ROM[3427] <= 12'h929; 
SIN_ROM[3428] <= 12'h92b; 
SIN_ROM[3429] <= 12'h92c; 
SIN_ROM[3430] <= 12'h92e; 
SIN_ROM[3431] <= 12'h930; 
SIN_ROM[3432] <= 12'h931; 
SIN_ROM[3433] <= 12'h933; 
SIN_ROM[3434] <= 12'h935; 
SIN_ROM[3435] <= 12'h936; 
SIN_ROM[3436] <= 12'h938; 
SIN_ROM[3437] <= 12'h93a; 
SIN_ROM[3438] <= 12'h93b; 
SIN_ROM[3439] <= 12'h93d; 
SIN_ROM[3440] <= 12'h93f; 
SIN_ROM[3441] <= 12'h940; 
SIN_ROM[3442] <= 12'h942; 
SIN_ROM[3443] <= 12'h944; 
SIN_ROM[3444] <= 12'h945; 
SIN_ROM[3445] <= 12'h947; 
SIN_ROM[3446] <= 12'h949; 
SIN_ROM[3447] <= 12'h94a; 
SIN_ROM[3448] <= 12'h94c; 
SIN_ROM[3449] <= 12'h94e; 
SIN_ROM[3450] <= 12'h950; 
SIN_ROM[3451] <= 12'h951; 
SIN_ROM[3452] <= 12'h953; 
SIN_ROM[3453] <= 12'h955; 
SIN_ROM[3454] <= 12'h957; 
SIN_ROM[3455] <= 12'h958; 
SIN_ROM[3456] <= 12'h95a; 
SIN_ROM[3457] <= 12'h95c; 
SIN_ROM[3458] <= 12'h95d; 
SIN_ROM[3459] <= 12'h95f; 
SIN_ROM[3460] <= 12'h961; 
SIN_ROM[3461] <= 12'h963; 
SIN_ROM[3462] <= 12'h965; 
SIN_ROM[3463] <= 12'h966; 
SIN_ROM[3464] <= 12'h968; 
SIN_ROM[3465] <= 12'h96a; 
SIN_ROM[3466] <= 12'h96c; 
SIN_ROM[3467] <= 12'h96d; 
SIN_ROM[3468] <= 12'h96f; 
SIN_ROM[3469] <= 12'h971; 
SIN_ROM[3470] <= 12'h973; 
SIN_ROM[3471] <= 12'h975; 
SIN_ROM[3472] <= 12'h976; 
SIN_ROM[3473] <= 12'h978; 
SIN_ROM[3474] <= 12'h97a; 
SIN_ROM[3475] <= 12'h97c; 
SIN_ROM[3476] <= 12'h97e; 
SIN_ROM[3477] <= 12'h97f; 
SIN_ROM[3478] <= 12'h981; 
SIN_ROM[3479] <= 12'h983; 
SIN_ROM[3480] <= 12'h985; 
SIN_ROM[3481] <= 12'h987; 
SIN_ROM[3482] <= 12'h989; 
SIN_ROM[3483] <= 12'h98b; 
SIN_ROM[3484] <= 12'h98c; 
SIN_ROM[3485] <= 12'h98e; 
SIN_ROM[3486] <= 12'h990; 
SIN_ROM[3487] <= 12'h992; 
SIN_ROM[3488] <= 12'h994; 
SIN_ROM[3489] <= 12'h996; 
SIN_ROM[3490] <= 12'h998; 
SIN_ROM[3491] <= 12'h999; 
SIN_ROM[3492] <= 12'h99b; 
SIN_ROM[3493] <= 12'h99d; 
SIN_ROM[3494] <= 12'h99f; 
SIN_ROM[3495] <= 12'h9a1; 
SIN_ROM[3496] <= 12'h9a3; 
SIN_ROM[3497] <= 12'h9a5; 
SIN_ROM[3498] <= 12'h9a7; 
SIN_ROM[3499] <= 12'h9a9; 
SIN_ROM[3500] <= 12'h9ab; 
SIN_ROM[3501] <= 12'h9ac; 
SIN_ROM[3502] <= 12'h9ae; 
SIN_ROM[3503] <= 12'h9b0; 
SIN_ROM[3504] <= 12'h9b2; 
SIN_ROM[3505] <= 12'h9b4; 
SIN_ROM[3506] <= 12'h9b6; 
SIN_ROM[3507] <= 12'h9b8; 
SIN_ROM[3508] <= 12'h9ba; 
SIN_ROM[3509] <= 12'h9bc; 
SIN_ROM[3510] <= 12'h9be; 
SIN_ROM[3511] <= 12'h9c0; 
SIN_ROM[3512] <= 12'h9c2; 
SIN_ROM[3513] <= 12'h9c4; 
SIN_ROM[3514] <= 12'h9c6; 
SIN_ROM[3515] <= 12'h9c8; 
SIN_ROM[3516] <= 12'h9ca; 
SIN_ROM[3517] <= 12'h9cc; 
SIN_ROM[3518] <= 12'h9ce; 
SIN_ROM[3519] <= 12'h9d0; 
SIN_ROM[3520] <= 12'h9d2; 
SIN_ROM[3521] <= 12'h9d4; 
SIN_ROM[3522] <= 12'h9d6; 
SIN_ROM[3523] <= 12'h9d8; 
SIN_ROM[3524] <= 12'h9da; 
SIN_ROM[3525] <= 12'h9dc; 
SIN_ROM[3526] <= 12'h9de; 
SIN_ROM[3527] <= 12'h9e0; 
SIN_ROM[3528] <= 12'h9e2; 
SIN_ROM[3529] <= 12'h9e4; 
SIN_ROM[3530] <= 12'h9e6; 
SIN_ROM[3531] <= 12'h9e8; 
SIN_ROM[3532] <= 12'h9ea; 
SIN_ROM[3533] <= 12'h9ec; 
SIN_ROM[3534] <= 12'h9ee; 
SIN_ROM[3535] <= 12'h9f0; 
SIN_ROM[3536] <= 12'h9f2; 
SIN_ROM[3537] <= 12'h9f4; 
SIN_ROM[3538] <= 12'h9f6; 
SIN_ROM[3539] <= 12'h9f8; 
SIN_ROM[3540] <= 12'h9fa; 
SIN_ROM[3541] <= 12'h9fc; 
SIN_ROM[3542] <= 12'h9fe; 
SIN_ROM[3543] <= 12'ha00; 
SIN_ROM[3544] <= 12'ha03; 
SIN_ROM[3545] <= 12'ha05; 
SIN_ROM[3546] <= 12'ha07; 
SIN_ROM[3547] <= 12'ha09; 
SIN_ROM[3548] <= 12'ha0b; 
SIN_ROM[3549] <= 12'ha0d; 
SIN_ROM[3550] <= 12'ha0f; 
SIN_ROM[3551] <= 12'ha11; 
SIN_ROM[3552] <= 12'ha13; 
SIN_ROM[3553] <= 12'ha15; 
SIN_ROM[3554] <= 12'ha17; 
SIN_ROM[3555] <= 12'ha1a; 
SIN_ROM[3556] <= 12'ha1c; 
SIN_ROM[3557] <= 12'ha1e; 
SIN_ROM[3558] <= 12'ha20; 
SIN_ROM[3559] <= 12'ha22; 
SIN_ROM[3560] <= 12'ha24; 
SIN_ROM[3561] <= 12'ha26; 
SIN_ROM[3562] <= 12'ha29; 
SIN_ROM[3563] <= 12'ha2b; 
SIN_ROM[3564] <= 12'ha2d; 
SIN_ROM[3565] <= 12'ha2f; 
SIN_ROM[3566] <= 12'ha31; 
SIN_ROM[3567] <= 12'ha33; 
SIN_ROM[3568] <= 12'ha35; 
SIN_ROM[3569] <= 12'ha38; 
SIN_ROM[3570] <= 12'ha3a; 
SIN_ROM[3571] <= 12'ha3c; 
SIN_ROM[3572] <= 12'ha3e; 
SIN_ROM[3573] <= 12'ha40; 
SIN_ROM[3574] <= 12'ha43; 
SIN_ROM[3575] <= 12'ha45; 
SIN_ROM[3576] <= 12'ha47; 
SIN_ROM[3577] <= 12'ha49; 
SIN_ROM[3578] <= 12'ha4b; 
SIN_ROM[3579] <= 12'ha4d; 
SIN_ROM[3580] <= 12'ha50; 
SIN_ROM[3581] <= 12'ha52; 
SIN_ROM[3582] <= 12'ha54; 
SIN_ROM[3583] <= 12'ha56; 
SIN_ROM[3584] <= 12'ha59; 
SIN_ROM[3585] <= 12'ha5b; 
SIN_ROM[3586] <= 12'ha5d; 
SIN_ROM[3587] <= 12'ha5f; 
SIN_ROM[3588] <= 12'ha61; 
SIN_ROM[3589] <= 12'ha64; 
SIN_ROM[3590] <= 12'ha66; 
SIN_ROM[3591] <= 12'ha68; 
SIN_ROM[3592] <= 12'ha6a; 
SIN_ROM[3593] <= 12'ha6d; 
SIN_ROM[3594] <= 12'ha6f; 
SIN_ROM[3595] <= 12'ha71; 
SIN_ROM[3596] <= 12'ha73; 
SIN_ROM[3597] <= 12'ha76; 
SIN_ROM[3598] <= 12'ha78; 
SIN_ROM[3599] <= 12'ha7a; 
SIN_ROM[3600] <= 12'ha7d; 
SIN_ROM[3601] <= 12'ha7f; 
SIN_ROM[3602] <= 12'ha81; 
SIN_ROM[3603] <= 12'ha83; 
SIN_ROM[3604] <= 12'ha86; 
SIN_ROM[3605] <= 12'ha88; 
SIN_ROM[3606] <= 12'ha8a; 
SIN_ROM[3607] <= 12'ha8d; 
SIN_ROM[3608] <= 12'ha8f; 
SIN_ROM[3609] <= 12'ha91; 
SIN_ROM[3610] <= 12'ha93; 
SIN_ROM[3611] <= 12'ha96; 
SIN_ROM[3612] <= 12'ha98; 
SIN_ROM[3613] <= 12'ha9a; 
SIN_ROM[3614] <= 12'ha9d; 
SIN_ROM[3615] <= 12'ha9f; 
SIN_ROM[3616] <= 12'haa1; 
SIN_ROM[3617] <= 12'haa4; 
SIN_ROM[3618] <= 12'haa6; 
SIN_ROM[3619] <= 12'haa8; 
SIN_ROM[3620] <= 12'haab; 
SIN_ROM[3621] <= 12'haad; 
SIN_ROM[3622] <= 12'haaf; 
SIN_ROM[3623] <= 12'hab2; 
SIN_ROM[3624] <= 12'hab4; 
SIN_ROM[3625] <= 12'hab6; 
SIN_ROM[3626] <= 12'hab9; 
SIN_ROM[3627] <= 12'habb; 
SIN_ROM[3628] <= 12'habd; 
SIN_ROM[3629] <= 12'hac0; 
SIN_ROM[3630] <= 12'hac2; 
SIN_ROM[3631] <= 12'hac5; 
SIN_ROM[3632] <= 12'hac7; 
SIN_ROM[3633] <= 12'hac9; 
SIN_ROM[3634] <= 12'hacc; 
SIN_ROM[3635] <= 12'hace; 
SIN_ROM[3636] <= 12'had0; 
SIN_ROM[3637] <= 12'had3; 
SIN_ROM[3638] <= 12'had5; 
SIN_ROM[3639] <= 12'had8; 
SIN_ROM[3640] <= 12'hada; 
SIN_ROM[3641] <= 12'hadc; 
SIN_ROM[3642] <= 12'hadf; 
SIN_ROM[3643] <= 12'hae1; 
SIN_ROM[3644] <= 12'hae4; 
SIN_ROM[3645] <= 12'hae6; 
SIN_ROM[3646] <= 12'hae9; 
SIN_ROM[3647] <= 12'haeb; 
SIN_ROM[3648] <= 12'haed; 
SIN_ROM[3649] <= 12'haf0; 
SIN_ROM[3650] <= 12'haf2; 
SIN_ROM[3651] <= 12'haf5; 
SIN_ROM[3652] <= 12'haf7; 
SIN_ROM[3653] <= 12'hafa; 
SIN_ROM[3654] <= 12'hafc; 
SIN_ROM[3655] <= 12'hafe; 
SIN_ROM[3656] <= 12'hb01; 
SIN_ROM[3657] <= 12'hb03; 
SIN_ROM[3658] <= 12'hb06; 
SIN_ROM[3659] <= 12'hb08; 
SIN_ROM[3660] <= 12'hb0b; 
SIN_ROM[3661] <= 12'hb0d; 
SIN_ROM[3662] <= 12'hb10; 
SIN_ROM[3663] <= 12'hb12; 
SIN_ROM[3664] <= 12'hb15; 
SIN_ROM[3665] <= 12'hb17; 
SIN_ROM[3666] <= 12'hb1a; 
SIN_ROM[3667] <= 12'hb1c; 
SIN_ROM[3668] <= 12'hb1f; 
SIN_ROM[3669] <= 12'hb21; 
SIN_ROM[3670] <= 12'hb24; 
SIN_ROM[3671] <= 12'hb26; 
SIN_ROM[3672] <= 12'hb29; 
SIN_ROM[3673] <= 12'hb2b; 
SIN_ROM[3674] <= 12'hb2e; 
SIN_ROM[3675] <= 12'hb30; 
SIN_ROM[3676] <= 12'hb33; 
SIN_ROM[3677] <= 12'hb35; 
SIN_ROM[3678] <= 12'hb38; 
SIN_ROM[3679] <= 12'hb3a; 
SIN_ROM[3680] <= 12'hb3d; 
SIN_ROM[3681] <= 12'hb3f; 
SIN_ROM[3682] <= 12'hb42; 
SIN_ROM[3683] <= 12'hb44; 
SIN_ROM[3684] <= 12'hb47; 
SIN_ROM[3685] <= 12'hb49; 
SIN_ROM[3686] <= 12'hb4c; 
SIN_ROM[3687] <= 12'hb4e; 
SIN_ROM[3688] <= 12'hb51; 
SIN_ROM[3689] <= 12'hb53; 
SIN_ROM[3690] <= 12'hb56; 
SIN_ROM[3691] <= 12'hb59; 
SIN_ROM[3692] <= 12'hb5b; 
SIN_ROM[3693] <= 12'hb5e; 
SIN_ROM[3694] <= 12'hb60; 
SIN_ROM[3695] <= 12'hb63; 
SIN_ROM[3696] <= 12'hb65; 
SIN_ROM[3697] <= 12'hb68; 
SIN_ROM[3698] <= 12'hb6a; 
SIN_ROM[3699] <= 12'hb6d; 
SIN_ROM[3700] <= 12'hb70; 
SIN_ROM[3701] <= 12'hb72; 
SIN_ROM[3702] <= 12'hb75; 
SIN_ROM[3703] <= 12'hb77; 
SIN_ROM[3704] <= 12'hb7a; 
SIN_ROM[3705] <= 12'hb7d; 
SIN_ROM[3706] <= 12'hb7f; 
SIN_ROM[3707] <= 12'hb82; 
SIN_ROM[3708] <= 12'hb84; 
SIN_ROM[3709] <= 12'hb87; 
SIN_ROM[3710] <= 12'hb8a; 
SIN_ROM[3711] <= 12'hb8c; 
SIN_ROM[3712] <= 12'hb8f; 
SIN_ROM[3713] <= 12'hb91; 
SIN_ROM[3714] <= 12'hb94; 
SIN_ROM[3715] <= 12'hb97; 
SIN_ROM[3716] <= 12'hb99; 
SIN_ROM[3717] <= 12'hb9c; 
SIN_ROM[3718] <= 12'hb9e; 
SIN_ROM[3719] <= 12'hba1; 
SIN_ROM[3720] <= 12'hba4; 
SIN_ROM[3721] <= 12'hba6; 
SIN_ROM[3722] <= 12'hba9; 
SIN_ROM[3723] <= 12'hbac; 
SIN_ROM[3724] <= 12'hbae; 
SIN_ROM[3725] <= 12'hbb1; 
SIN_ROM[3726] <= 12'hbb4; 
SIN_ROM[3727] <= 12'hbb6; 
SIN_ROM[3728] <= 12'hbb9; 
SIN_ROM[3729] <= 12'hbbc; 
SIN_ROM[3730] <= 12'hbbe; 
SIN_ROM[3731] <= 12'hbc1; 
SIN_ROM[3732] <= 12'hbc3; 
SIN_ROM[3733] <= 12'hbc6; 
SIN_ROM[3734] <= 12'hbc9; 
SIN_ROM[3735] <= 12'hbcb; 
SIN_ROM[3736] <= 12'hbce; 
SIN_ROM[3737] <= 12'hbd1; 
SIN_ROM[3738] <= 12'hbd4; 
SIN_ROM[3739] <= 12'hbd6; 
SIN_ROM[3740] <= 12'hbd9; 
SIN_ROM[3741] <= 12'hbdc; 
SIN_ROM[3742] <= 12'hbde; 
SIN_ROM[3743] <= 12'hbe1; 
SIN_ROM[3744] <= 12'hbe4; 
SIN_ROM[3745] <= 12'hbe6; 
SIN_ROM[3746] <= 12'hbe9; 
SIN_ROM[3747] <= 12'hbec; 
SIN_ROM[3748] <= 12'hbee; 
SIN_ROM[3749] <= 12'hbf1; 
SIN_ROM[3750] <= 12'hbf4; 
SIN_ROM[3751] <= 12'hbf7; 
SIN_ROM[3752] <= 12'hbf9; 
SIN_ROM[3753] <= 12'hbfc; 
SIN_ROM[3754] <= 12'hbff; 
SIN_ROM[3755] <= 12'hc01; 
SIN_ROM[3756] <= 12'hc04; 
SIN_ROM[3757] <= 12'hc07; 
SIN_ROM[3758] <= 12'hc0a; 
SIN_ROM[3759] <= 12'hc0c; 
SIN_ROM[3760] <= 12'hc0f; 
SIN_ROM[3761] <= 12'hc12; 
SIN_ROM[3762] <= 12'hc15; 
SIN_ROM[3763] <= 12'hc17; 
SIN_ROM[3764] <= 12'hc1a; 
SIN_ROM[3765] <= 12'hc1d; 
SIN_ROM[3766] <= 12'hc1f; 
SIN_ROM[3767] <= 12'hc22; 
SIN_ROM[3768] <= 12'hc25; 
SIN_ROM[3769] <= 12'hc28; 
SIN_ROM[3770] <= 12'hc2a; 
SIN_ROM[3771] <= 12'hc2d; 
SIN_ROM[3772] <= 12'hc30; 
SIN_ROM[3773] <= 12'hc33; 
SIN_ROM[3774] <= 12'hc36; 
SIN_ROM[3775] <= 12'hc38; 
SIN_ROM[3776] <= 12'hc3b; 
SIN_ROM[3777] <= 12'hc3e; 
SIN_ROM[3778] <= 12'hc41; 
SIN_ROM[3779] <= 12'hc43; 
SIN_ROM[3780] <= 12'hc46; 
SIN_ROM[3781] <= 12'hc49; 
SIN_ROM[3782] <= 12'hc4c; 
SIN_ROM[3783] <= 12'hc4e; 
SIN_ROM[3784] <= 12'hc51; 
SIN_ROM[3785] <= 12'hc54; 
SIN_ROM[3786] <= 12'hc57; 
SIN_ROM[3787] <= 12'hc5a; 
SIN_ROM[3788] <= 12'hc5c; 
SIN_ROM[3789] <= 12'hc5f; 
SIN_ROM[3790] <= 12'hc62; 
SIN_ROM[3791] <= 12'hc65; 
SIN_ROM[3792] <= 12'hc68; 
SIN_ROM[3793] <= 12'hc6a; 
SIN_ROM[3794] <= 12'hc6d; 
SIN_ROM[3795] <= 12'hc70; 
SIN_ROM[3796] <= 12'hc73; 
SIN_ROM[3797] <= 12'hc76; 
SIN_ROM[3798] <= 12'hc79; 
SIN_ROM[3799] <= 12'hc7b; 
SIN_ROM[3800] <= 12'hc7e; 
SIN_ROM[3801] <= 12'hc81; 
SIN_ROM[3802] <= 12'hc84; 
SIN_ROM[3803] <= 12'hc87; 
SIN_ROM[3804] <= 12'hc89; 
SIN_ROM[3805] <= 12'hc8c; 
SIN_ROM[3806] <= 12'hc8f; 
SIN_ROM[3807] <= 12'hc92; 
SIN_ROM[3808] <= 12'hc95; 
SIN_ROM[3809] <= 12'hc98; 
SIN_ROM[3810] <= 12'hc9a; 
SIN_ROM[3811] <= 12'hc9d; 
SIN_ROM[3812] <= 12'hca0; 
SIN_ROM[3813] <= 12'hca3; 
SIN_ROM[3814] <= 12'hca6; 
SIN_ROM[3815] <= 12'hca9; 
SIN_ROM[3816] <= 12'hcac; 
SIN_ROM[3817] <= 12'hcae; 
SIN_ROM[3818] <= 12'hcb1; 
SIN_ROM[3819] <= 12'hcb4; 
SIN_ROM[3820] <= 12'hcb7; 
SIN_ROM[3821] <= 12'hcba; 
SIN_ROM[3822] <= 12'hcbd; 
SIN_ROM[3823] <= 12'hcc0; 
SIN_ROM[3824] <= 12'hcc2; 
SIN_ROM[3825] <= 12'hcc5; 
SIN_ROM[3826] <= 12'hcc8; 
SIN_ROM[3827] <= 12'hccb; 
SIN_ROM[3828] <= 12'hcce; 
SIN_ROM[3829] <= 12'hcd1; 
SIN_ROM[3830] <= 12'hcd4; 
SIN_ROM[3831] <= 12'hcd7; 
SIN_ROM[3832] <= 12'hcd9; 
SIN_ROM[3833] <= 12'hcdc; 
SIN_ROM[3834] <= 12'hcdf; 
SIN_ROM[3835] <= 12'hce2; 
SIN_ROM[3836] <= 12'hce5; 
SIN_ROM[3837] <= 12'hce8; 
SIN_ROM[3838] <= 12'hceb; 
SIN_ROM[3839] <= 12'hcee; 
SIN_ROM[3840] <= 12'hcf1; 
SIN_ROM[3841] <= 12'hcf4; 
SIN_ROM[3842] <= 12'hcf6; 
SIN_ROM[3843] <= 12'hcf9; 
SIN_ROM[3844] <= 12'hcfc; 
SIN_ROM[3845] <= 12'hcff; 
SIN_ROM[3846] <= 12'hd02; 
SIN_ROM[3847] <= 12'hd05; 
SIN_ROM[3848] <= 12'hd08; 
SIN_ROM[3849] <= 12'hd0b; 
SIN_ROM[3850] <= 12'hd0e; 
SIN_ROM[3851] <= 12'hd11; 
SIN_ROM[3852] <= 12'hd14; 
SIN_ROM[3853] <= 12'hd17; 
SIN_ROM[3854] <= 12'hd19; 
SIN_ROM[3855] <= 12'hd1c; 
SIN_ROM[3856] <= 12'hd1f; 
SIN_ROM[3857] <= 12'hd22; 
SIN_ROM[3858] <= 12'hd25; 
SIN_ROM[3859] <= 12'hd28; 
SIN_ROM[3860] <= 12'hd2b; 
SIN_ROM[3861] <= 12'hd2e; 
SIN_ROM[3862] <= 12'hd31; 
SIN_ROM[3863] <= 12'hd34; 
SIN_ROM[3864] <= 12'hd37; 
SIN_ROM[3865] <= 12'hd3a; 
SIN_ROM[3866] <= 12'hd3d; 
SIN_ROM[3867] <= 12'hd40; 
SIN_ROM[3868] <= 12'hd43; 
SIN_ROM[3869] <= 12'hd46; 
SIN_ROM[3870] <= 12'hd48; 
SIN_ROM[3871] <= 12'hd4b; 
SIN_ROM[3872] <= 12'hd4e; 
SIN_ROM[3873] <= 12'hd51; 
SIN_ROM[3874] <= 12'hd54; 
SIN_ROM[3875] <= 12'hd57; 
SIN_ROM[3876] <= 12'hd5a; 
SIN_ROM[3877] <= 12'hd5d; 
SIN_ROM[3878] <= 12'hd60; 
SIN_ROM[3879] <= 12'hd63; 
SIN_ROM[3880] <= 12'hd66; 
SIN_ROM[3881] <= 12'hd69; 
SIN_ROM[3882] <= 12'hd6c; 
SIN_ROM[3883] <= 12'hd6f; 
SIN_ROM[3884] <= 12'hd72; 
SIN_ROM[3885] <= 12'hd75; 
SIN_ROM[3886] <= 12'hd78; 
SIN_ROM[3887] <= 12'hd7b; 
SIN_ROM[3888] <= 12'hd7e; 
SIN_ROM[3889] <= 12'hd81; 
SIN_ROM[3890] <= 12'hd84; 
SIN_ROM[3891] <= 12'hd87; 
SIN_ROM[3892] <= 12'hd8a; 
SIN_ROM[3893] <= 12'hd8d; 
SIN_ROM[3894] <= 12'hd90; 
SIN_ROM[3895] <= 12'hd93; 
SIN_ROM[3896] <= 12'hd96; 
SIN_ROM[3897] <= 12'hd99; 
SIN_ROM[3898] <= 12'hd9c; 
SIN_ROM[3899] <= 12'hd9f; 
SIN_ROM[3900] <= 12'hda2; 
SIN_ROM[3901] <= 12'hda5; 
SIN_ROM[3902] <= 12'hda8; 
SIN_ROM[3903] <= 12'hdab; 
SIN_ROM[3904] <= 12'hdae; 
SIN_ROM[3905] <= 12'hdb1; 
SIN_ROM[3906] <= 12'hdb4; 
SIN_ROM[3907] <= 12'hdb7; 
SIN_ROM[3908] <= 12'hdba; 
SIN_ROM[3909] <= 12'hdbd; 
SIN_ROM[3910] <= 12'hdc0; 
SIN_ROM[3911] <= 12'hdc3; 
SIN_ROM[3912] <= 12'hdc6; 
SIN_ROM[3913] <= 12'hdc9; 
SIN_ROM[3914] <= 12'hdcc; 
SIN_ROM[3915] <= 12'hdcf; 
SIN_ROM[3916] <= 12'hdd2; 
SIN_ROM[3917] <= 12'hdd5; 
SIN_ROM[3918] <= 12'hdd8; 
SIN_ROM[3919] <= 12'hddb; 
SIN_ROM[3920] <= 12'hdde; 
SIN_ROM[3921] <= 12'hde1; 
SIN_ROM[3922] <= 12'hde4; 
SIN_ROM[3923] <= 12'hde7; 
SIN_ROM[3924] <= 12'hdea; 
SIN_ROM[3925] <= 12'hded; 
SIN_ROM[3926] <= 12'hdf0; 
SIN_ROM[3927] <= 12'hdf3; 
SIN_ROM[3928] <= 12'hdf6; 
SIN_ROM[3929] <= 12'hdf9; 
SIN_ROM[3930] <= 12'hdfc; 
SIN_ROM[3931] <= 12'hdff; 
SIN_ROM[3932] <= 12'he02; 
SIN_ROM[3933] <= 12'he05; 
SIN_ROM[3934] <= 12'he09; 
SIN_ROM[3935] <= 12'he0c; 
SIN_ROM[3936] <= 12'he0f; 
SIN_ROM[3937] <= 12'he12; 
SIN_ROM[3938] <= 12'he15; 
SIN_ROM[3939] <= 12'he18; 
SIN_ROM[3940] <= 12'he1b; 
SIN_ROM[3941] <= 12'he1e; 
SIN_ROM[3942] <= 12'he21; 
SIN_ROM[3943] <= 12'he24; 
SIN_ROM[3944] <= 12'he27; 
SIN_ROM[3945] <= 12'he2a; 
SIN_ROM[3946] <= 12'he2d; 
SIN_ROM[3947] <= 12'he30; 
SIN_ROM[3948] <= 12'he33; 
SIN_ROM[3949] <= 12'he36; 
SIN_ROM[3950] <= 12'he39; 
SIN_ROM[3951] <= 12'he3c; 
SIN_ROM[3952] <= 12'he3f; 
SIN_ROM[3953] <= 12'he43; 
SIN_ROM[3954] <= 12'he46; 
SIN_ROM[3955] <= 12'he49; 
SIN_ROM[3956] <= 12'he4c; 
SIN_ROM[3957] <= 12'he4f; 
SIN_ROM[3958] <= 12'he52; 
SIN_ROM[3959] <= 12'he55; 
SIN_ROM[3960] <= 12'he58; 
SIN_ROM[3961] <= 12'he5b; 
SIN_ROM[3962] <= 12'he5e; 
SIN_ROM[3963] <= 12'he61; 
SIN_ROM[3964] <= 12'he64; 
SIN_ROM[3965] <= 12'he67; 
SIN_ROM[3966] <= 12'he6a; 
SIN_ROM[3967] <= 12'he6e; 
SIN_ROM[3968] <= 12'he71; 
SIN_ROM[3969] <= 12'he74; 
SIN_ROM[3970] <= 12'he77; 
SIN_ROM[3971] <= 12'he7a; 
SIN_ROM[3972] <= 12'he7d; 
SIN_ROM[3973] <= 12'he80; 
SIN_ROM[3974] <= 12'he83; 
SIN_ROM[3975] <= 12'he86; 
SIN_ROM[3976] <= 12'he89; 
SIN_ROM[3977] <= 12'he8c; 
SIN_ROM[3978] <= 12'he8f; 
SIN_ROM[3979] <= 12'he93; 
SIN_ROM[3980] <= 12'he96; 
SIN_ROM[3981] <= 12'he99; 
SIN_ROM[3982] <= 12'he9c; 
SIN_ROM[3983] <= 12'he9f; 
SIN_ROM[3984] <= 12'hea2; 
SIN_ROM[3985] <= 12'hea5; 
SIN_ROM[3986] <= 12'hea8; 
SIN_ROM[3987] <= 12'heab; 
SIN_ROM[3988] <= 12'heae; 
SIN_ROM[3989] <= 12'heb2; 
SIN_ROM[3990] <= 12'heb5; 
SIN_ROM[3991] <= 12'heb8; 
SIN_ROM[3992] <= 12'hebb; 
SIN_ROM[3993] <= 12'hebe; 
SIN_ROM[3994] <= 12'hec1; 
SIN_ROM[3995] <= 12'hec4; 
SIN_ROM[3996] <= 12'hec7; 
SIN_ROM[3997] <= 12'heca; 
SIN_ROM[3998] <= 12'hecd; 
SIN_ROM[3999] <= 12'hed1; 
SIN_ROM[4000] <= 12'hed4; 
SIN_ROM[4001] <= 12'hed7; 
SIN_ROM[4002] <= 12'heda; 
SIN_ROM[4003] <= 12'hedd; 
SIN_ROM[4004] <= 12'hee0; 
SIN_ROM[4005] <= 12'hee3; 
SIN_ROM[4006] <= 12'hee6; 
SIN_ROM[4007] <= 12'hee9; 
SIN_ROM[4008] <= 12'heed; 
SIN_ROM[4009] <= 12'hef0; 
SIN_ROM[4010] <= 12'hef3; 
SIN_ROM[4011] <= 12'hef6; 
SIN_ROM[4012] <= 12'hef9; 
SIN_ROM[4013] <= 12'hefc; 
SIN_ROM[4014] <= 12'heff; 
SIN_ROM[4015] <= 12'hf02; 
SIN_ROM[4016] <= 12'hf05; 
SIN_ROM[4017] <= 12'hf09; 
SIN_ROM[4018] <= 12'hf0c; 
SIN_ROM[4019] <= 12'hf0f; 
SIN_ROM[4020] <= 12'hf12; 
SIN_ROM[4021] <= 12'hf15; 
SIN_ROM[4022] <= 12'hf18; 
SIN_ROM[4023] <= 12'hf1b; 
SIN_ROM[4024] <= 12'hf1e; 
SIN_ROM[4025] <= 12'hf21; 
SIN_ROM[4026] <= 12'hf25; 
SIN_ROM[4027] <= 12'hf28; 
SIN_ROM[4028] <= 12'hf2b; 
SIN_ROM[4029] <= 12'hf2e; 
SIN_ROM[4030] <= 12'hf31; 
SIN_ROM[4031] <= 12'hf34; 
SIN_ROM[4032] <= 12'hf37; 
SIN_ROM[4033] <= 12'hf3a; 
SIN_ROM[4034] <= 12'hf3e; 
SIN_ROM[4035] <= 12'hf41; 
SIN_ROM[4036] <= 12'hf44; 
SIN_ROM[4037] <= 12'hf47; 
SIN_ROM[4038] <= 12'hf4a; 
SIN_ROM[4039] <= 12'hf4d; 
SIN_ROM[4040] <= 12'hf50; 
SIN_ROM[4041] <= 12'hf54; 
SIN_ROM[4042] <= 12'hf57; 
SIN_ROM[4043] <= 12'hf5a; 
SIN_ROM[4044] <= 12'hf5d; 
SIN_ROM[4045] <= 12'hf60; 
SIN_ROM[4046] <= 12'hf63; 
SIN_ROM[4047] <= 12'hf66; 
SIN_ROM[4048] <= 12'hf69; 
SIN_ROM[4049] <= 12'hf6d; 
SIN_ROM[4050] <= 12'hf70; 
SIN_ROM[4051] <= 12'hf73; 
SIN_ROM[4052] <= 12'hf76; 
SIN_ROM[4053] <= 12'hf79; 
SIN_ROM[4054] <= 12'hf7c; 
SIN_ROM[4055] <= 12'hf7f; 
SIN_ROM[4056] <= 12'hf82; 
SIN_ROM[4057] <= 12'hf86; 
SIN_ROM[4058] <= 12'hf89; 
SIN_ROM[4059] <= 12'hf8c; 
SIN_ROM[4060] <= 12'hf8f; 
SIN_ROM[4061] <= 12'hf92; 
SIN_ROM[4062] <= 12'hf95; 
SIN_ROM[4063] <= 12'hf98; 
SIN_ROM[4064] <= 12'hf9c; 
SIN_ROM[4065] <= 12'hf9f; 
SIN_ROM[4066] <= 12'hfa2; 
SIN_ROM[4067] <= 12'hfa5; 
SIN_ROM[4068] <= 12'hfa8; 
SIN_ROM[4069] <= 12'hfab; 
SIN_ROM[4070] <= 12'hfae; 
SIN_ROM[4071] <= 12'hfb2; 
SIN_ROM[4072] <= 12'hfb5; 
SIN_ROM[4073] <= 12'hfb8; 
SIN_ROM[4074] <= 12'hfbb; 
SIN_ROM[4075] <= 12'hfbe; 
SIN_ROM[4076] <= 12'hfc1; 
SIN_ROM[4077] <= 12'hfc4; 
SIN_ROM[4078] <= 12'hfc7; 
SIN_ROM[4079] <= 12'hfcb; 
SIN_ROM[4080] <= 12'hfce; 
SIN_ROM[4081] <= 12'hfd1; 
SIN_ROM[4082] <= 12'hfd4; 
SIN_ROM[4083] <= 12'hfd7; 
SIN_ROM[4084] <= 12'hfda; 
SIN_ROM[4085] <= 12'hfdd; 
SIN_ROM[4086] <= 12'hfe1; 
SIN_ROM[4087] <= 12'hfe4; 
SIN_ROM[4088] <= 12'hfe7; 
SIN_ROM[4089] <= 12'hfea; 
SIN_ROM[4090] <= 12'hfed; 
SIN_ROM[4091] <= 12'hff0; 
SIN_ROM[4092] <= 12'hff3; 
SIN_ROM[4093] <= 12'hff7; 
SIN_ROM[4094] <= 12'hffa; 
SIN_ROM[4095] <= 12'hffd; 


COS_ROM[0] <= 12'h7ff; 
COS_ROM[1] <= 12'h7ff; 
COS_ROM[2] <= 12'h7ff; 
COS_ROM[3] <= 12'h7ff; 
COS_ROM[4] <= 12'h7ff; 
COS_ROM[5] <= 12'h7ff; 
COS_ROM[6] <= 12'h7ff; 
COS_ROM[7] <= 12'h7ff; 
COS_ROM[8] <= 12'h7ff; 
COS_ROM[9] <= 12'h7ff; 
COS_ROM[10] <= 12'h7ff; 
COS_ROM[11] <= 12'h7ff; 
COS_ROM[12] <= 12'h7ff; 
COS_ROM[13] <= 12'h7ff; 
COS_ROM[14] <= 12'h7ff; 
COS_ROM[15] <= 12'h7fe; 
COS_ROM[16] <= 12'h7fe; 
COS_ROM[17] <= 12'h7fe; 
COS_ROM[18] <= 12'h7fe; 
COS_ROM[19] <= 12'h7fe; 
COS_ROM[20] <= 12'h7fe; 
COS_ROM[21] <= 12'h7fe; 
COS_ROM[22] <= 12'h7fe; 
COS_ROM[23] <= 12'h7fe; 
COS_ROM[24] <= 12'h7fe; 
COS_ROM[25] <= 12'h7fd; 
COS_ROM[26] <= 12'h7fd; 
COS_ROM[27] <= 12'h7fd; 
COS_ROM[28] <= 12'h7fd; 
COS_ROM[29] <= 12'h7fd; 
COS_ROM[30] <= 12'h7fd; 
COS_ROM[31] <= 12'h7fd; 
COS_ROM[32] <= 12'h7fd; 
COS_ROM[33] <= 12'h7fc; 
COS_ROM[34] <= 12'h7fc; 
COS_ROM[35] <= 12'h7fc; 
COS_ROM[36] <= 12'h7fc; 
COS_ROM[37] <= 12'h7fc; 
COS_ROM[38] <= 12'h7fc; 
COS_ROM[39] <= 12'h7fb; 
COS_ROM[40] <= 12'h7fb; 
COS_ROM[41] <= 12'h7fb; 
COS_ROM[42] <= 12'h7fb; 
COS_ROM[43] <= 12'h7fb; 
COS_ROM[44] <= 12'h7fa; 
COS_ROM[45] <= 12'h7fa; 
COS_ROM[46] <= 12'h7fa; 
COS_ROM[47] <= 12'h7fa; 
COS_ROM[48] <= 12'h7f9; 
COS_ROM[49] <= 12'h7f9; 
COS_ROM[50] <= 12'h7f9; 
COS_ROM[51] <= 12'h7f9; 
COS_ROM[52] <= 12'h7f8; 
COS_ROM[53] <= 12'h7f8; 
COS_ROM[54] <= 12'h7f8; 
COS_ROM[55] <= 12'h7f8; 
COS_ROM[56] <= 12'h7f7; 
COS_ROM[57] <= 12'h7f7; 
COS_ROM[58] <= 12'h7f7; 
COS_ROM[59] <= 12'h7f7; 
COS_ROM[60] <= 12'h7f6; 
COS_ROM[61] <= 12'h7f6; 
COS_ROM[62] <= 12'h7f6; 
COS_ROM[63] <= 12'h7f5; 
COS_ROM[64] <= 12'h7f5; 
COS_ROM[65] <= 12'h7f5; 
COS_ROM[66] <= 12'h7f5; 
COS_ROM[67] <= 12'h7f4; 
COS_ROM[68] <= 12'h7f4; 
COS_ROM[69] <= 12'h7f4; 
COS_ROM[70] <= 12'h7f3; 
COS_ROM[71] <= 12'h7f3; 
COS_ROM[72] <= 12'h7f3; 
COS_ROM[73] <= 12'h7f2; 
COS_ROM[74] <= 12'h7f2; 
COS_ROM[75] <= 12'h7f1; 
COS_ROM[76] <= 12'h7f1; 
COS_ROM[77] <= 12'h7f1; 
COS_ROM[78] <= 12'h7f0; 
COS_ROM[79] <= 12'h7f0; 
COS_ROM[80] <= 12'h7f0; 
COS_ROM[81] <= 12'h7ef; 
COS_ROM[82] <= 12'h7ef; 
COS_ROM[83] <= 12'h7ee; 
COS_ROM[84] <= 12'h7ee; 
COS_ROM[85] <= 12'h7ee; 
COS_ROM[86] <= 12'h7ed; 
COS_ROM[87] <= 12'h7ed; 
COS_ROM[88] <= 12'h7ec; 
COS_ROM[89] <= 12'h7ec; 
COS_ROM[90] <= 12'h7ec; 
COS_ROM[91] <= 12'h7eb; 
COS_ROM[92] <= 12'h7eb; 
COS_ROM[93] <= 12'h7ea; 
COS_ROM[94] <= 12'h7ea; 
COS_ROM[95] <= 12'h7e9; 
COS_ROM[96] <= 12'h7e9; 
COS_ROM[97] <= 12'h7e8; 
COS_ROM[98] <= 12'h7e8; 
COS_ROM[99] <= 12'h7e7; 
COS_ROM[100] <= 12'h7e7; 
COS_ROM[101] <= 12'h7e6; 
COS_ROM[102] <= 12'h7e6; 
COS_ROM[103] <= 12'h7e6; 
COS_ROM[104] <= 12'h7e5; 
COS_ROM[105] <= 12'h7e5; 
COS_ROM[106] <= 12'h7e4; 
COS_ROM[107] <= 12'h7e3; 
COS_ROM[108] <= 12'h7e3; 
COS_ROM[109] <= 12'h7e2; 
COS_ROM[110] <= 12'h7e2; 
COS_ROM[111] <= 12'h7e1; 
COS_ROM[112] <= 12'h7e1; 
COS_ROM[113] <= 12'h7e0; 
COS_ROM[114] <= 12'h7e0; 
COS_ROM[115] <= 12'h7df; 
COS_ROM[116] <= 12'h7df; 
COS_ROM[117] <= 12'h7de; 
COS_ROM[118] <= 12'h7de; 
COS_ROM[119] <= 12'h7dd; 
COS_ROM[120] <= 12'h7dc; 
COS_ROM[121] <= 12'h7dc; 
COS_ROM[122] <= 12'h7db; 
COS_ROM[123] <= 12'h7db; 
COS_ROM[124] <= 12'h7da; 
COS_ROM[125] <= 12'h7d9; 
COS_ROM[126] <= 12'h7d9; 
COS_ROM[127] <= 12'h7d8; 
COS_ROM[128] <= 12'h7d8; 
COS_ROM[129] <= 12'h7d7; 
COS_ROM[130] <= 12'h7d6; 
COS_ROM[131] <= 12'h7d6; 
COS_ROM[132] <= 12'h7d5; 
COS_ROM[133] <= 12'h7d5; 
COS_ROM[134] <= 12'h7d4; 
COS_ROM[135] <= 12'h7d3; 
COS_ROM[136] <= 12'h7d3; 
COS_ROM[137] <= 12'h7d2; 
COS_ROM[138] <= 12'h7d1; 
COS_ROM[139] <= 12'h7d1; 
COS_ROM[140] <= 12'h7d0; 
COS_ROM[141] <= 12'h7cf; 
COS_ROM[142] <= 12'h7cf; 
COS_ROM[143] <= 12'h7ce; 
COS_ROM[144] <= 12'h7cd; 
COS_ROM[145] <= 12'h7cd; 
COS_ROM[146] <= 12'h7cc; 
COS_ROM[147] <= 12'h7cb; 
COS_ROM[148] <= 12'h7ca; 
COS_ROM[149] <= 12'h7ca; 
COS_ROM[150] <= 12'h7c9; 
COS_ROM[151] <= 12'h7c8; 
COS_ROM[152] <= 12'h7c8; 
COS_ROM[153] <= 12'h7c7; 
COS_ROM[154] <= 12'h7c6; 
COS_ROM[155] <= 12'h7c5; 
COS_ROM[156] <= 12'h7c5; 
COS_ROM[157] <= 12'h7c4; 
COS_ROM[158] <= 12'h7c3; 
COS_ROM[159] <= 12'h7c2; 
COS_ROM[160] <= 12'h7c2; 
COS_ROM[161] <= 12'h7c1; 
COS_ROM[162] <= 12'h7c0; 
COS_ROM[163] <= 12'h7bf; 
COS_ROM[164] <= 12'h7bf; 
COS_ROM[165] <= 12'h7be; 
COS_ROM[166] <= 12'h7bd; 
COS_ROM[167] <= 12'h7bc; 
COS_ROM[168] <= 12'h7bb; 
COS_ROM[169] <= 12'h7bb; 
COS_ROM[170] <= 12'h7ba; 
COS_ROM[171] <= 12'h7b9; 
COS_ROM[172] <= 12'h7b8; 
COS_ROM[173] <= 12'h7b7; 
COS_ROM[174] <= 12'h7b7; 
COS_ROM[175] <= 12'h7b6; 
COS_ROM[176] <= 12'h7b5; 
COS_ROM[177] <= 12'h7b4; 
COS_ROM[178] <= 12'h7b3; 
COS_ROM[179] <= 12'h7b2; 
COS_ROM[180] <= 12'h7b1; 
COS_ROM[181] <= 12'h7b1; 
COS_ROM[182] <= 12'h7b0; 
COS_ROM[183] <= 12'h7af; 
COS_ROM[184] <= 12'h7ae; 
COS_ROM[185] <= 12'h7ad; 
COS_ROM[186] <= 12'h7ac; 
COS_ROM[187] <= 12'h7ab; 
COS_ROM[188] <= 12'h7aa; 
COS_ROM[189] <= 12'h7aa; 
COS_ROM[190] <= 12'h7a9; 
COS_ROM[191] <= 12'h7a8; 
COS_ROM[192] <= 12'h7a7; 
COS_ROM[193] <= 12'h7a6; 
COS_ROM[194] <= 12'h7a5; 
COS_ROM[195] <= 12'h7a4; 
COS_ROM[196] <= 12'h7a3; 
COS_ROM[197] <= 12'h7a2; 
COS_ROM[198] <= 12'h7a1; 
COS_ROM[199] <= 12'h7a0; 
COS_ROM[200] <= 12'h79f; 
COS_ROM[201] <= 12'h79e; 
COS_ROM[202] <= 12'h79e; 
COS_ROM[203] <= 12'h79d; 
COS_ROM[204] <= 12'h79c; 
COS_ROM[205] <= 12'h79b; 
COS_ROM[206] <= 12'h79a; 
COS_ROM[207] <= 12'h799; 
COS_ROM[208] <= 12'h798; 
COS_ROM[209] <= 12'h797; 
COS_ROM[210] <= 12'h796; 
COS_ROM[211] <= 12'h795; 
COS_ROM[212] <= 12'h794; 
COS_ROM[213] <= 12'h793; 
COS_ROM[214] <= 12'h792; 
COS_ROM[215] <= 12'h791; 
COS_ROM[216] <= 12'h790; 
COS_ROM[217] <= 12'h78f; 
COS_ROM[218] <= 12'h78e; 
COS_ROM[219] <= 12'h78d; 
COS_ROM[220] <= 12'h78c; 
COS_ROM[221] <= 12'h78a; 
COS_ROM[222] <= 12'h789; 
COS_ROM[223] <= 12'h788; 
COS_ROM[224] <= 12'h787; 
COS_ROM[225] <= 12'h786; 
COS_ROM[226] <= 12'h785; 
COS_ROM[227] <= 12'h784; 
COS_ROM[228] <= 12'h783; 
COS_ROM[229] <= 12'h782; 
COS_ROM[230] <= 12'h781; 
COS_ROM[231] <= 12'h780; 
COS_ROM[232] <= 12'h77f; 
COS_ROM[233] <= 12'h77e; 
COS_ROM[234] <= 12'h77d; 
COS_ROM[235] <= 12'h77b; 
COS_ROM[236] <= 12'h77a; 
COS_ROM[237] <= 12'h779; 
COS_ROM[238] <= 12'h778; 
COS_ROM[239] <= 12'h777; 
COS_ROM[240] <= 12'h776; 
COS_ROM[241] <= 12'h775; 
COS_ROM[242] <= 12'h774; 
COS_ROM[243] <= 12'h772; 
COS_ROM[244] <= 12'h771; 
COS_ROM[245] <= 12'h770; 
COS_ROM[246] <= 12'h76f; 
COS_ROM[247] <= 12'h76e; 
COS_ROM[248] <= 12'h76d; 
COS_ROM[249] <= 12'h76b; 
COS_ROM[250] <= 12'h76a; 
COS_ROM[251] <= 12'h769; 
COS_ROM[252] <= 12'h768; 
COS_ROM[253] <= 12'h767; 
COS_ROM[254] <= 12'h766; 
COS_ROM[255] <= 12'h764; 
COS_ROM[256] <= 12'h763; 
COS_ROM[257] <= 12'h762; 
COS_ROM[258] <= 12'h761; 
COS_ROM[259] <= 12'h760; 
COS_ROM[260] <= 12'h75e; 
COS_ROM[261] <= 12'h75d; 
COS_ROM[262] <= 12'h75c; 
COS_ROM[263] <= 12'h75b; 
COS_ROM[264] <= 12'h759; 
COS_ROM[265] <= 12'h758; 
COS_ROM[266] <= 12'h757; 
COS_ROM[267] <= 12'h756; 
COS_ROM[268] <= 12'h754; 
COS_ROM[269] <= 12'h753; 
COS_ROM[270] <= 12'h752; 
COS_ROM[271] <= 12'h751; 
COS_ROM[272] <= 12'h74f; 
COS_ROM[273] <= 12'h74e; 
COS_ROM[274] <= 12'h74d; 
COS_ROM[275] <= 12'h74c; 
COS_ROM[276] <= 12'h74a; 
COS_ROM[277] <= 12'h749; 
COS_ROM[278] <= 12'h748; 
COS_ROM[279] <= 12'h746; 
COS_ROM[280] <= 12'h745; 
COS_ROM[281] <= 12'h744; 
COS_ROM[282] <= 12'h742; 
COS_ROM[283] <= 12'h741; 
COS_ROM[284] <= 12'h740; 
COS_ROM[285] <= 12'h73e; 
COS_ROM[286] <= 12'h73d; 
COS_ROM[287] <= 12'h73c; 
COS_ROM[288] <= 12'h73a; 
COS_ROM[289] <= 12'h739; 
COS_ROM[290] <= 12'h738; 
COS_ROM[291] <= 12'h736; 
COS_ROM[292] <= 12'h735; 
COS_ROM[293] <= 12'h734; 
COS_ROM[294] <= 12'h732; 
COS_ROM[295] <= 12'h731; 
COS_ROM[296] <= 12'h730; 
COS_ROM[297] <= 12'h72e; 
COS_ROM[298] <= 12'h72d; 
COS_ROM[299] <= 12'h72b; 
COS_ROM[300] <= 12'h72a; 
COS_ROM[301] <= 12'h729; 
COS_ROM[302] <= 12'h727; 
COS_ROM[303] <= 12'h726; 
COS_ROM[304] <= 12'h724; 
COS_ROM[305] <= 12'h723; 
COS_ROM[306] <= 12'h722; 
COS_ROM[307] <= 12'h720; 
COS_ROM[308] <= 12'h71f; 
COS_ROM[309] <= 12'h71d; 
COS_ROM[310] <= 12'h71c; 
COS_ROM[311] <= 12'h71a; 
COS_ROM[312] <= 12'h719; 
COS_ROM[313] <= 12'h718; 
COS_ROM[314] <= 12'h716; 
COS_ROM[315] <= 12'h715; 
COS_ROM[316] <= 12'h713; 
COS_ROM[317] <= 12'h712; 
COS_ROM[318] <= 12'h710; 
COS_ROM[319] <= 12'h70f; 
COS_ROM[320] <= 12'h70d; 
COS_ROM[321] <= 12'h70c; 
COS_ROM[322] <= 12'h70a; 
COS_ROM[323] <= 12'h709; 
COS_ROM[324] <= 12'h707; 
COS_ROM[325] <= 12'h706; 
COS_ROM[326] <= 12'h704; 
COS_ROM[327] <= 12'h703; 
COS_ROM[328] <= 12'h701; 
COS_ROM[329] <= 12'h700; 
COS_ROM[330] <= 12'h6fe; 
COS_ROM[331] <= 12'h6fd; 
COS_ROM[332] <= 12'h6fb; 
COS_ROM[333] <= 12'h6fa; 
COS_ROM[334] <= 12'h6f8; 
COS_ROM[335] <= 12'h6f7; 
COS_ROM[336] <= 12'h6f5; 
COS_ROM[337] <= 12'h6f4; 
COS_ROM[338] <= 12'h6f2; 
COS_ROM[339] <= 12'h6f0; 
COS_ROM[340] <= 12'h6ef; 
COS_ROM[341] <= 12'h6ed; 
COS_ROM[342] <= 12'h6ec; 
COS_ROM[343] <= 12'h6ea; 
COS_ROM[344] <= 12'h6e9; 
COS_ROM[345] <= 12'h6e7; 
COS_ROM[346] <= 12'h6e5; 
COS_ROM[347] <= 12'h6e4; 
COS_ROM[348] <= 12'h6e2; 
COS_ROM[349] <= 12'h6e1; 
COS_ROM[350] <= 12'h6df; 
COS_ROM[351] <= 12'h6dd; 
COS_ROM[352] <= 12'h6dc; 
COS_ROM[353] <= 12'h6da; 
COS_ROM[354] <= 12'h6d9; 
COS_ROM[355] <= 12'h6d7; 
COS_ROM[356] <= 12'h6d5; 
COS_ROM[357] <= 12'h6d4; 
COS_ROM[358] <= 12'h6d2; 
COS_ROM[359] <= 12'h6d0; 
COS_ROM[360] <= 12'h6cf; 
COS_ROM[361] <= 12'h6cd; 
COS_ROM[362] <= 12'h6cb; 
COS_ROM[363] <= 12'h6ca; 
COS_ROM[364] <= 12'h6c8; 
COS_ROM[365] <= 12'h6c6; 
COS_ROM[366] <= 12'h6c5; 
COS_ROM[367] <= 12'h6c3; 
COS_ROM[368] <= 12'h6c1; 
COS_ROM[369] <= 12'h6c0; 
COS_ROM[370] <= 12'h6be; 
COS_ROM[371] <= 12'h6bc; 
COS_ROM[372] <= 12'h6bb; 
COS_ROM[373] <= 12'h6b9; 
COS_ROM[374] <= 12'h6b7; 
COS_ROM[375] <= 12'h6b6; 
COS_ROM[376] <= 12'h6b4; 
COS_ROM[377] <= 12'h6b2; 
COS_ROM[378] <= 12'h6b0; 
COS_ROM[379] <= 12'h6af; 
COS_ROM[380] <= 12'h6ad; 
COS_ROM[381] <= 12'h6ab; 
COS_ROM[382] <= 12'h6a9; 
COS_ROM[383] <= 12'h6a8; 
COS_ROM[384] <= 12'h6a6; 
COS_ROM[385] <= 12'h6a4; 
COS_ROM[386] <= 12'h6a3; 
COS_ROM[387] <= 12'h6a1; 
COS_ROM[388] <= 12'h69f; 
COS_ROM[389] <= 12'h69d; 
COS_ROM[390] <= 12'h69b; 
COS_ROM[391] <= 12'h69a; 
COS_ROM[392] <= 12'h698; 
COS_ROM[393] <= 12'h696; 
COS_ROM[394] <= 12'h694; 
COS_ROM[395] <= 12'h693; 
COS_ROM[396] <= 12'h691; 
COS_ROM[397] <= 12'h68f; 
COS_ROM[398] <= 12'h68d; 
COS_ROM[399] <= 12'h68b; 
COS_ROM[400] <= 12'h68a; 
COS_ROM[401] <= 12'h688; 
COS_ROM[402] <= 12'h686; 
COS_ROM[403] <= 12'h684; 
COS_ROM[404] <= 12'h682; 
COS_ROM[405] <= 12'h681; 
COS_ROM[406] <= 12'h67f; 
COS_ROM[407] <= 12'h67d; 
COS_ROM[408] <= 12'h67b; 
COS_ROM[409] <= 12'h679; 
COS_ROM[410] <= 12'h677; 
COS_ROM[411] <= 12'h675; 
COS_ROM[412] <= 12'h674; 
COS_ROM[413] <= 12'h672; 
COS_ROM[414] <= 12'h670; 
COS_ROM[415] <= 12'h66e; 
COS_ROM[416] <= 12'h66c; 
COS_ROM[417] <= 12'h66a; 
COS_ROM[418] <= 12'h668; 
COS_ROM[419] <= 12'h667; 
COS_ROM[420] <= 12'h665; 
COS_ROM[421] <= 12'h663; 
COS_ROM[422] <= 12'h661; 
COS_ROM[423] <= 12'h65f; 
COS_ROM[424] <= 12'h65d; 
COS_ROM[425] <= 12'h65b; 
COS_ROM[426] <= 12'h659; 
COS_ROM[427] <= 12'h657; 
COS_ROM[428] <= 12'h655; 
COS_ROM[429] <= 12'h654; 
COS_ROM[430] <= 12'h652; 
COS_ROM[431] <= 12'h650; 
COS_ROM[432] <= 12'h64e; 
COS_ROM[433] <= 12'h64c; 
COS_ROM[434] <= 12'h64a; 
COS_ROM[435] <= 12'h648; 
COS_ROM[436] <= 12'h646; 
COS_ROM[437] <= 12'h644; 
COS_ROM[438] <= 12'h642; 
COS_ROM[439] <= 12'h640; 
COS_ROM[440] <= 12'h63e; 
COS_ROM[441] <= 12'h63c; 
COS_ROM[442] <= 12'h63a; 
COS_ROM[443] <= 12'h638; 
COS_ROM[444] <= 12'h636; 
COS_ROM[445] <= 12'h634; 
COS_ROM[446] <= 12'h632; 
COS_ROM[447] <= 12'h630; 
COS_ROM[448] <= 12'h62e; 
COS_ROM[449] <= 12'h62c; 
COS_ROM[450] <= 12'h62a; 
COS_ROM[451] <= 12'h628; 
COS_ROM[452] <= 12'h626; 
COS_ROM[453] <= 12'h624; 
COS_ROM[454] <= 12'h622; 
COS_ROM[455] <= 12'h620; 
COS_ROM[456] <= 12'h61e; 
COS_ROM[457] <= 12'h61c; 
COS_ROM[458] <= 12'h61a; 
COS_ROM[459] <= 12'h618; 
COS_ROM[460] <= 12'h616; 
COS_ROM[461] <= 12'h614; 
COS_ROM[462] <= 12'h612; 
COS_ROM[463] <= 12'h610; 
COS_ROM[464] <= 12'h60e; 
COS_ROM[465] <= 12'h60c; 
COS_ROM[466] <= 12'h60a; 
COS_ROM[467] <= 12'h608; 
COS_ROM[468] <= 12'h606; 
COS_ROM[469] <= 12'h604; 
COS_ROM[470] <= 12'h602; 
COS_ROM[471] <= 12'h600; 
COS_ROM[472] <= 12'h5fd; 
COS_ROM[473] <= 12'h5fb; 
COS_ROM[474] <= 12'h5f9; 
COS_ROM[475] <= 12'h5f7; 
COS_ROM[476] <= 12'h5f5; 
COS_ROM[477] <= 12'h5f3; 
COS_ROM[478] <= 12'h5f1; 
COS_ROM[479] <= 12'h5ef; 
COS_ROM[480] <= 12'h5ed; 
COS_ROM[481] <= 12'h5eb; 
COS_ROM[482] <= 12'h5e9; 
COS_ROM[483] <= 12'h5e6; 
COS_ROM[484] <= 12'h5e4; 
COS_ROM[485] <= 12'h5e2; 
COS_ROM[486] <= 12'h5e0; 
COS_ROM[487] <= 12'h5de; 
COS_ROM[488] <= 12'h5dc; 
COS_ROM[489] <= 12'h5da; 
COS_ROM[490] <= 12'h5d7; 
COS_ROM[491] <= 12'h5d5; 
COS_ROM[492] <= 12'h5d3; 
COS_ROM[493] <= 12'h5d1; 
COS_ROM[494] <= 12'h5cf; 
COS_ROM[495] <= 12'h5cd; 
COS_ROM[496] <= 12'h5cb; 
COS_ROM[497] <= 12'h5c8; 
COS_ROM[498] <= 12'h5c6; 
COS_ROM[499] <= 12'h5c4; 
COS_ROM[500] <= 12'h5c2; 
COS_ROM[501] <= 12'h5c0; 
COS_ROM[502] <= 12'h5bd; 
COS_ROM[503] <= 12'h5bb; 
COS_ROM[504] <= 12'h5b9; 
COS_ROM[505] <= 12'h5b7; 
COS_ROM[506] <= 12'h5b5; 
COS_ROM[507] <= 12'h5b3; 
COS_ROM[508] <= 12'h5b0; 
COS_ROM[509] <= 12'h5ae; 
COS_ROM[510] <= 12'h5ac; 
COS_ROM[511] <= 12'h5aa; 
COS_ROM[512] <= 12'h5a7; 
COS_ROM[513] <= 12'h5a5; 
COS_ROM[514] <= 12'h5a3; 
COS_ROM[515] <= 12'h5a1; 
COS_ROM[516] <= 12'h59f; 
COS_ROM[517] <= 12'h59c; 
COS_ROM[518] <= 12'h59a; 
COS_ROM[519] <= 12'h598; 
COS_ROM[520] <= 12'h596; 
COS_ROM[521] <= 12'h593; 
COS_ROM[522] <= 12'h591; 
COS_ROM[523] <= 12'h58f; 
COS_ROM[524] <= 12'h58d; 
COS_ROM[525] <= 12'h58a; 
COS_ROM[526] <= 12'h588; 
COS_ROM[527] <= 12'h586; 
COS_ROM[528] <= 12'h583; 
COS_ROM[529] <= 12'h581; 
COS_ROM[530] <= 12'h57f; 
COS_ROM[531] <= 12'h57d; 
COS_ROM[532] <= 12'h57a; 
COS_ROM[533] <= 12'h578; 
COS_ROM[534] <= 12'h576; 
COS_ROM[535] <= 12'h573; 
COS_ROM[536] <= 12'h571; 
COS_ROM[537] <= 12'h56f; 
COS_ROM[538] <= 12'h56d; 
COS_ROM[539] <= 12'h56a; 
COS_ROM[540] <= 12'h568; 
COS_ROM[541] <= 12'h566; 
COS_ROM[542] <= 12'h563; 
COS_ROM[543] <= 12'h561; 
COS_ROM[544] <= 12'h55f; 
COS_ROM[545] <= 12'h55c; 
COS_ROM[546] <= 12'h55a; 
COS_ROM[547] <= 12'h558; 
COS_ROM[548] <= 12'h555; 
COS_ROM[549] <= 12'h553; 
COS_ROM[550] <= 12'h551; 
COS_ROM[551] <= 12'h54e; 
COS_ROM[552] <= 12'h54c; 
COS_ROM[553] <= 12'h54a; 
COS_ROM[554] <= 12'h547; 
COS_ROM[555] <= 12'h545; 
COS_ROM[556] <= 12'h543; 
COS_ROM[557] <= 12'h540; 
COS_ROM[558] <= 12'h53e; 
COS_ROM[559] <= 12'h53b; 
COS_ROM[560] <= 12'h539; 
COS_ROM[561] <= 12'h537; 
COS_ROM[562] <= 12'h534; 
COS_ROM[563] <= 12'h532; 
COS_ROM[564] <= 12'h530; 
COS_ROM[565] <= 12'h52d; 
COS_ROM[566] <= 12'h52b; 
COS_ROM[567] <= 12'h528; 
COS_ROM[568] <= 12'h526; 
COS_ROM[569] <= 12'h524; 
COS_ROM[570] <= 12'h521; 
COS_ROM[571] <= 12'h51f; 
COS_ROM[572] <= 12'h51c; 
COS_ROM[573] <= 12'h51a; 
COS_ROM[574] <= 12'h517; 
COS_ROM[575] <= 12'h515; 
COS_ROM[576] <= 12'h513; 
COS_ROM[577] <= 12'h510; 
COS_ROM[578] <= 12'h50e; 
COS_ROM[579] <= 12'h50b; 
COS_ROM[580] <= 12'h509; 
COS_ROM[581] <= 12'h506; 
COS_ROM[582] <= 12'h504; 
COS_ROM[583] <= 12'h502; 
COS_ROM[584] <= 12'h4ff; 
COS_ROM[585] <= 12'h4fd; 
COS_ROM[586] <= 12'h4fa; 
COS_ROM[587] <= 12'h4f8; 
COS_ROM[588] <= 12'h4f5; 
COS_ROM[589] <= 12'h4f3; 
COS_ROM[590] <= 12'h4f0; 
COS_ROM[591] <= 12'h4ee; 
COS_ROM[592] <= 12'h4eb; 
COS_ROM[593] <= 12'h4e9; 
COS_ROM[594] <= 12'h4e6; 
COS_ROM[595] <= 12'h4e4; 
COS_ROM[596] <= 12'h4e1; 
COS_ROM[597] <= 12'h4df; 
COS_ROM[598] <= 12'h4dc; 
COS_ROM[599] <= 12'h4da; 
COS_ROM[600] <= 12'h4d7; 
COS_ROM[601] <= 12'h4d5; 
COS_ROM[602] <= 12'h4d2; 
COS_ROM[603] <= 12'h4d0; 
COS_ROM[604] <= 12'h4cd; 
COS_ROM[605] <= 12'h4cb; 
COS_ROM[606] <= 12'h4c8; 
COS_ROM[607] <= 12'h4c6; 
COS_ROM[608] <= 12'h4c3; 
COS_ROM[609] <= 12'h4c1; 
COS_ROM[610] <= 12'h4be; 
COS_ROM[611] <= 12'h4bc; 
COS_ROM[612] <= 12'h4b9; 
COS_ROM[613] <= 12'h4b7; 
COS_ROM[614] <= 12'h4b4; 
COS_ROM[615] <= 12'h4b2; 
COS_ROM[616] <= 12'h4af; 
COS_ROM[617] <= 12'h4ad; 
COS_ROM[618] <= 12'h4aa; 
COS_ROM[619] <= 12'h4a7; 
COS_ROM[620] <= 12'h4a5; 
COS_ROM[621] <= 12'h4a2; 
COS_ROM[622] <= 12'h4a0; 
COS_ROM[623] <= 12'h49d; 
COS_ROM[624] <= 12'h49b; 
COS_ROM[625] <= 12'h498; 
COS_ROM[626] <= 12'h496; 
COS_ROM[627] <= 12'h493; 
COS_ROM[628] <= 12'h490; 
COS_ROM[629] <= 12'h48e; 
COS_ROM[630] <= 12'h48b; 
COS_ROM[631] <= 12'h489; 
COS_ROM[632] <= 12'h486; 
COS_ROM[633] <= 12'h483; 
COS_ROM[634] <= 12'h481; 
COS_ROM[635] <= 12'h47e; 
COS_ROM[636] <= 12'h47c; 
COS_ROM[637] <= 12'h479; 
COS_ROM[638] <= 12'h476; 
COS_ROM[639] <= 12'h474; 
COS_ROM[640] <= 12'h471; 
COS_ROM[641] <= 12'h46f; 
COS_ROM[642] <= 12'h46c; 
COS_ROM[643] <= 12'h469; 
COS_ROM[644] <= 12'h467; 
COS_ROM[645] <= 12'h464; 
COS_ROM[646] <= 12'h462; 
COS_ROM[647] <= 12'h45f; 
COS_ROM[648] <= 12'h45c; 
COS_ROM[649] <= 12'h45a; 
COS_ROM[650] <= 12'h457; 
COS_ROM[651] <= 12'h454; 
COS_ROM[652] <= 12'h452; 
COS_ROM[653] <= 12'h44f; 
COS_ROM[654] <= 12'h44c; 
COS_ROM[655] <= 12'h44a; 
COS_ROM[656] <= 12'h447; 
COS_ROM[657] <= 12'h444; 
COS_ROM[658] <= 12'h442; 
COS_ROM[659] <= 12'h43f; 
COS_ROM[660] <= 12'h43d; 
COS_ROM[661] <= 12'h43a; 
COS_ROM[662] <= 12'h437; 
COS_ROM[663] <= 12'h435; 
COS_ROM[664] <= 12'h432; 
COS_ROM[665] <= 12'h42f; 
COS_ROM[666] <= 12'h42c; 
COS_ROM[667] <= 12'h42a; 
COS_ROM[668] <= 12'h427; 
COS_ROM[669] <= 12'h424; 
COS_ROM[670] <= 12'h422; 
COS_ROM[671] <= 12'h41f; 
COS_ROM[672] <= 12'h41c; 
COS_ROM[673] <= 12'h41a; 
COS_ROM[674] <= 12'h417; 
COS_ROM[675] <= 12'h414; 
COS_ROM[676] <= 12'h412; 
COS_ROM[677] <= 12'h40f; 
COS_ROM[678] <= 12'h40c; 
COS_ROM[679] <= 12'h409; 
COS_ROM[680] <= 12'h407; 
COS_ROM[681] <= 12'h404; 
COS_ROM[682] <= 12'h401; 
COS_ROM[683] <= 12'h3ff; 
COS_ROM[684] <= 12'h3fc; 
COS_ROM[685] <= 12'h3f9; 
COS_ROM[686] <= 12'h3f6; 
COS_ROM[687] <= 12'h3f4; 
COS_ROM[688] <= 12'h3f1; 
COS_ROM[689] <= 12'h3ee; 
COS_ROM[690] <= 12'h3eb; 
COS_ROM[691] <= 12'h3e9; 
COS_ROM[692] <= 12'h3e6; 
COS_ROM[693] <= 12'h3e3; 
COS_ROM[694] <= 12'h3e1; 
COS_ROM[695] <= 12'h3de; 
COS_ROM[696] <= 12'h3db; 
COS_ROM[697] <= 12'h3d8; 
COS_ROM[698] <= 12'h3d6; 
COS_ROM[699] <= 12'h3d3; 
COS_ROM[700] <= 12'h3d0; 
COS_ROM[701] <= 12'h3cd; 
COS_ROM[702] <= 12'h3ca; 
COS_ROM[703] <= 12'h3c8; 
COS_ROM[704] <= 12'h3c5; 
COS_ROM[705] <= 12'h3c2; 
COS_ROM[706] <= 12'h3bf; 
COS_ROM[707] <= 12'h3bd; 
COS_ROM[708] <= 12'h3ba; 
COS_ROM[709] <= 12'h3b7; 
COS_ROM[710] <= 12'h3b4; 
COS_ROM[711] <= 12'h3b2; 
COS_ROM[712] <= 12'h3af; 
COS_ROM[713] <= 12'h3ac; 
COS_ROM[714] <= 12'h3a9; 
COS_ROM[715] <= 12'h3a6; 
COS_ROM[716] <= 12'h3a4; 
COS_ROM[717] <= 12'h3a1; 
COS_ROM[718] <= 12'h39e; 
COS_ROM[719] <= 12'h39b; 
COS_ROM[720] <= 12'h398; 
COS_ROM[721] <= 12'h396; 
COS_ROM[722] <= 12'h393; 
COS_ROM[723] <= 12'h390; 
COS_ROM[724] <= 12'h38d; 
COS_ROM[725] <= 12'h38a; 
COS_ROM[726] <= 12'h387; 
COS_ROM[727] <= 12'h385; 
COS_ROM[728] <= 12'h382; 
COS_ROM[729] <= 12'h37f; 
COS_ROM[730] <= 12'h37c; 
COS_ROM[731] <= 12'h379; 
COS_ROM[732] <= 12'h377; 
COS_ROM[733] <= 12'h374; 
COS_ROM[734] <= 12'h371; 
COS_ROM[735] <= 12'h36e; 
COS_ROM[736] <= 12'h36b; 
COS_ROM[737] <= 12'h368; 
COS_ROM[738] <= 12'h366; 
COS_ROM[739] <= 12'h363; 
COS_ROM[740] <= 12'h360; 
COS_ROM[741] <= 12'h35d; 
COS_ROM[742] <= 12'h35a; 
COS_ROM[743] <= 12'h357; 
COS_ROM[744] <= 12'h354; 
COS_ROM[745] <= 12'h352; 
COS_ROM[746] <= 12'h34f; 
COS_ROM[747] <= 12'h34c; 
COS_ROM[748] <= 12'h349; 
COS_ROM[749] <= 12'h346; 
COS_ROM[750] <= 12'h343; 
COS_ROM[751] <= 12'h340; 
COS_ROM[752] <= 12'h33e; 
COS_ROM[753] <= 12'h33b; 
COS_ROM[754] <= 12'h338; 
COS_ROM[755] <= 12'h335; 
COS_ROM[756] <= 12'h332; 
COS_ROM[757] <= 12'h32f; 
COS_ROM[758] <= 12'h32c; 
COS_ROM[759] <= 12'h329; 
COS_ROM[760] <= 12'h327; 
COS_ROM[761] <= 12'h324; 
COS_ROM[762] <= 12'h321; 
COS_ROM[763] <= 12'h31e; 
COS_ROM[764] <= 12'h31b; 
COS_ROM[765] <= 12'h318; 
COS_ROM[766] <= 12'h315; 
COS_ROM[767] <= 12'h312; 
COS_ROM[768] <= 12'h30f; 
COS_ROM[769] <= 12'h30c; 
COS_ROM[770] <= 12'h30a; 
COS_ROM[771] <= 12'h307; 
COS_ROM[772] <= 12'h304; 
COS_ROM[773] <= 12'h301; 
COS_ROM[774] <= 12'h2fe; 
COS_ROM[775] <= 12'h2fb; 
COS_ROM[776] <= 12'h2f8; 
COS_ROM[777] <= 12'h2f5; 
COS_ROM[778] <= 12'h2f2; 
COS_ROM[779] <= 12'h2ef; 
COS_ROM[780] <= 12'h2ec; 
COS_ROM[781] <= 12'h2e9; 
COS_ROM[782] <= 12'h2e7; 
COS_ROM[783] <= 12'h2e4; 
COS_ROM[784] <= 12'h2e1; 
COS_ROM[785] <= 12'h2de; 
COS_ROM[786] <= 12'h2db; 
COS_ROM[787] <= 12'h2d8; 
COS_ROM[788] <= 12'h2d5; 
COS_ROM[789] <= 12'h2d2; 
COS_ROM[790] <= 12'h2cf; 
COS_ROM[791] <= 12'h2cc; 
COS_ROM[792] <= 12'h2c9; 
COS_ROM[793] <= 12'h2c6; 
COS_ROM[794] <= 12'h2c3; 
COS_ROM[795] <= 12'h2c0; 
COS_ROM[796] <= 12'h2bd; 
COS_ROM[797] <= 12'h2ba; 
COS_ROM[798] <= 12'h2b8; 
COS_ROM[799] <= 12'h2b5; 
COS_ROM[800] <= 12'h2b2; 
COS_ROM[801] <= 12'h2af; 
COS_ROM[802] <= 12'h2ac; 
COS_ROM[803] <= 12'h2a9; 
COS_ROM[804] <= 12'h2a6; 
COS_ROM[805] <= 12'h2a3; 
COS_ROM[806] <= 12'h2a0; 
COS_ROM[807] <= 12'h29d; 
COS_ROM[808] <= 12'h29a; 
COS_ROM[809] <= 12'h297; 
COS_ROM[810] <= 12'h294; 
COS_ROM[811] <= 12'h291; 
COS_ROM[812] <= 12'h28e; 
COS_ROM[813] <= 12'h28b; 
COS_ROM[814] <= 12'h288; 
COS_ROM[815] <= 12'h285; 
COS_ROM[816] <= 12'h282; 
COS_ROM[817] <= 12'h27f; 
COS_ROM[818] <= 12'h27c; 
COS_ROM[819] <= 12'h279; 
COS_ROM[820] <= 12'h276; 
COS_ROM[821] <= 12'h273; 
COS_ROM[822] <= 12'h270; 
COS_ROM[823] <= 12'h26d; 
COS_ROM[824] <= 12'h26a; 
COS_ROM[825] <= 12'h267; 
COS_ROM[826] <= 12'h264; 
COS_ROM[827] <= 12'h261; 
COS_ROM[828] <= 12'h25e; 
COS_ROM[829] <= 12'h25b; 
COS_ROM[830] <= 12'h258; 
COS_ROM[831] <= 12'h255; 
COS_ROM[832] <= 12'h252; 
COS_ROM[833] <= 12'h24f; 
COS_ROM[834] <= 12'h24c; 
COS_ROM[835] <= 12'h249; 
COS_ROM[836] <= 12'h246; 
COS_ROM[837] <= 12'h243; 
COS_ROM[838] <= 12'h240; 
COS_ROM[839] <= 12'h23d; 
COS_ROM[840] <= 12'h23a; 
COS_ROM[841] <= 12'h237; 
COS_ROM[842] <= 12'h234; 
COS_ROM[843] <= 12'h231; 
COS_ROM[844] <= 12'h22e; 
COS_ROM[845] <= 12'h22b; 
COS_ROM[846] <= 12'h228; 
COS_ROM[847] <= 12'h225; 
COS_ROM[848] <= 12'h222; 
COS_ROM[849] <= 12'h21f; 
COS_ROM[850] <= 12'h21c; 
COS_ROM[851] <= 12'h219; 
COS_ROM[852] <= 12'h216; 
COS_ROM[853] <= 12'h213; 
COS_ROM[854] <= 12'h210; 
COS_ROM[855] <= 12'h20d; 
COS_ROM[856] <= 12'h20a; 
COS_ROM[857] <= 12'h207; 
COS_ROM[858] <= 12'h204; 
COS_ROM[859] <= 12'h201; 
COS_ROM[860] <= 12'h1fe; 
COS_ROM[861] <= 12'h1fb; 
COS_ROM[862] <= 12'h1f7; 
COS_ROM[863] <= 12'h1f4; 
COS_ROM[864] <= 12'h1f1; 
COS_ROM[865] <= 12'h1ee; 
COS_ROM[866] <= 12'h1eb; 
COS_ROM[867] <= 12'h1e8; 
COS_ROM[868] <= 12'h1e5; 
COS_ROM[869] <= 12'h1e2; 
COS_ROM[870] <= 12'h1df; 
COS_ROM[871] <= 12'h1dc; 
COS_ROM[872] <= 12'h1d9; 
COS_ROM[873] <= 12'h1d6; 
COS_ROM[874] <= 12'h1d3; 
COS_ROM[875] <= 12'h1d0; 
COS_ROM[876] <= 12'h1cd; 
COS_ROM[877] <= 12'h1ca; 
COS_ROM[878] <= 12'h1c7; 
COS_ROM[879] <= 12'h1c4; 
COS_ROM[880] <= 12'h1c1; 
COS_ROM[881] <= 12'h1bd; 
COS_ROM[882] <= 12'h1ba; 
COS_ROM[883] <= 12'h1b7; 
COS_ROM[884] <= 12'h1b4; 
COS_ROM[885] <= 12'h1b1; 
COS_ROM[886] <= 12'h1ae; 
COS_ROM[887] <= 12'h1ab; 
COS_ROM[888] <= 12'h1a8; 
COS_ROM[889] <= 12'h1a5; 
COS_ROM[890] <= 12'h1a2; 
COS_ROM[891] <= 12'h19f; 
COS_ROM[892] <= 12'h19c; 
COS_ROM[893] <= 12'h199; 
COS_ROM[894] <= 12'h196; 
COS_ROM[895] <= 12'h192; 
COS_ROM[896] <= 12'h18f; 
COS_ROM[897] <= 12'h18c; 
COS_ROM[898] <= 12'h189; 
COS_ROM[899] <= 12'h186; 
COS_ROM[900] <= 12'h183; 
COS_ROM[901] <= 12'h180; 
COS_ROM[902] <= 12'h17d; 
COS_ROM[903] <= 12'h17a; 
COS_ROM[904] <= 12'h177; 
COS_ROM[905] <= 12'h174; 
COS_ROM[906] <= 12'h171; 
COS_ROM[907] <= 12'h16d; 
COS_ROM[908] <= 12'h16a; 
COS_ROM[909] <= 12'h167; 
COS_ROM[910] <= 12'h164; 
COS_ROM[911] <= 12'h161; 
COS_ROM[912] <= 12'h15e; 
COS_ROM[913] <= 12'h15b; 
COS_ROM[914] <= 12'h158; 
COS_ROM[915] <= 12'h155; 
COS_ROM[916] <= 12'h152; 
COS_ROM[917] <= 12'h14e; 
COS_ROM[918] <= 12'h14b; 
COS_ROM[919] <= 12'h148; 
COS_ROM[920] <= 12'h145; 
COS_ROM[921] <= 12'h142; 
COS_ROM[922] <= 12'h13f; 
COS_ROM[923] <= 12'h13c; 
COS_ROM[924] <= 12'h139; 
COS_ROM[925] <= 12'h136; 
COS_ROM[926] <= 12'h133; 
COS_ROM[927] <= 12'h12f; 
COS_ROM[928] <= 12'h12c; 
COS_ROM[929] <= 12'h129; 
COS_ROM[930] <= 12'h126; 
COS_ROM[931] <= 12'h123; 
COS_ROM[932] <= 12'h120; 
COS_ROM[933] <= 12'h11d; 
COS_ROM[934] <= 12'h11a; 
COS_ROM[935] <= 12'h117; 
COS_ROM[936] <= 12'h113; 
COS_ROM[937] <= 12'h110; 
COS_ROM[938] <= 12'h10d; 
COS_ROM[939] <= 12'h10a; 
COS_ROM[940] <= 12'h107; 
COS_ROM[941] <= 12'h104; 
COS_ROM[942] <= 12'h101; 
COS_ROM[943] <= 12'h0fe; 
COS_ROM[944] <= 12'h0fb; 
COS_ROM[945] <= 12'h0f7; 
COS_ROM[946] <= 12'h0f4; 
COS_ROM[947] <= 12'h0f1; 
COS_ROM[948] <= 12'h0ee; 
COS_ROM[949] <= 12'h0eb; 
COS_ROM[950] <= 12'h0e8; 
COS_ROM[951] <= 12'h0e5; 
COS_ROM[952] <= 12'h0e2; 
COS_ROM[953] <= 12'h0df; 
COS_ROM[954] <= 12'h0db; 
COS_ROM[955] <= 12'h0d8; 
COS_ROM[956] <= 12'h0d5; 
COS_ROM[957] <= 12'h0d2; 
COS_ROM[958] <= 12'h0cf; 
COS_ROM[959] <= 12'h0cc; 
COS_ROM[960] <= 12'h0c9; 
COS_ROM[961] <= 12'h0c6; 
COS_ROM[962] <= 12'h0c2; 
COS_ROM[963] <= 12'h0bf; 
COS_ROM[964] <= 12'h0bc; 
COS_ROM[965] <= 12'h0b9; 
COS_ROM[966] <= 12'h0b6; 
COS_ROM[967] <= 12'h0b3; 
COS_ROM[968] <= 12'h0b0; 
COS_ROM[969] <= 12'h0ac; 
COS_ROM[970] <= 12'h0a9; 
COS_ROM[971] <= 12'h0a6; 
COS_ROM[972] <= 12'h0a3; 
COS_ROM[973] <= 12'h0a0; 
COS_ROM[974] <= 12'h09d; 
COS_ROM[975] <= 12'h09a; 
COS_ROM[976] <= 12'h097; 
COS_ROM[977] <= 12'h093; 
COS_ROM[978] <= 12'h090; 
COS_ROM[979] <= 12'h08d; 
COS_ROM[980] <= 12'h08a; 
COS_ROM[981] <= 12'h087; 
COS_ROM[982] <= 12'h084; 
COS_ROM[983] <= 12'h081; 
COS_ROM[984] <= 12'h07e; 
COS_ROM[985] <= 12'h07a; 
COS_ROM[986] <= 12'h077; 
COS_ROM[987] <= 12'h074; 
COS_ROM[988] <= 12'h071; 
COS_ROM[989] <= 12'h06e; 
COS_ROM[990] <= 12'h06b; 
COS_ROM[991] <= 12'h068; 
COS_ROM[992] <= 12'h064; 
COS_ROM[993] <= 12'h061; 
COS_ROM[994] <= 12'h05e; 
COS_ROM[995] <= 12'h05b; 
COS_ROM[996] <= 12'h058; 
COS_ROM[997] <= 12'h055; 
COS_ROM[998] <= 12'h052; 
COS_ROM[999] <= 12'h04e; 
COS_ROM[1000] <= 12'h04b; 
COS_ROM[1001] <= 12'h048; 
COS_ROM[1002] <= 12'h045; 
COS_ROM[1003] <= 12'h042; 
COS_ROM[1004] <= 12'h03f; 
COS_ROM[1005] <= 12'h03c; 
COS_ROM[1006] <= 12'h039; 
COS_ROM[1007] <= 12'h035; 
COS_ROM[1008] <= 12'h032; 
COS_ROM[1009] <= 12'h02f; 
COS_ROM[1010] <= 12'h02c; 
COS_ROM[1011] <= 12'h029; 
COS_ROM[1012] <= 12'h026; 
COS_ROM[1013] <= 12'h023; 
COS_ROM[1014] <= 12'h01f; 
COS_ROM[1015] <= 12'h01c; 
COS_ROM[1016] <= 12'h019; 
COS_ROM[1017] <= 12'h016; 
COS_ROM[1018] <= 12'h013; 
COS_ROM[1019] <= 12'h010; 
COS_ROM[1020] <= 12'h00d; 
COS_ROM[1021] <= 12'h009; 
COS_ROM[1022] <= 12'h006; 
COS_ROM[1023] <= 12'h003; 
COS_ROM[1024] <= 12'h000; 
COS_ROM[1025] <= 12'hffd; 
COS_ROM[1026] <= 12'hffa; 
COS_ROM[1027] <= 12'hff7; 
COS_ROM[1028] <= 12'hff3; 
COS_ROM[1029] <= 12'hff0; 
COS_ROM[1030] <= 12'hfed; 
COS_ROM[1031] <= 12'hfea; 
COS_ROM[1032] <= 12'hfe7; 
COS_ROM[1033] <= 12'hfe4; 
COS_ROM[1034] <= 12'hfe1; 
COS_ROM[1035] <= 12'hfdd; 
COS_ROM[1036] <= 12'hfda; 
COS_ROM[1037] <= 12'hfd7; 
COS_ROM[1038] <= 12'hfd4; 
COS_ROM[1039] <= 12'hfd1; 
COS_ROM[1040] <= 12'hfce; 
COS_ROM[1041] <= 12'hfcb; 
COS_ROM[1042] <= 12'hfc7; 
COS_ROM[1043] <= 12'hfc4; 
COS_ROM[1044] <= 12'hfc1; 
COS_ROM[1045] <= 12'hfbe; 
COS_ROM[1046] <= 12'hfbb; 
COS_ROM[1047] <= 12'hfb8; 
COS_ROM[1048] <= 12'hfb5; 
COS_ROM[1049] <= 12'hfb2; 
COS_ROM[1050] <= 12'hfae; 
COS_ROM[1051] <= 12'hfab; 
COS_ROM[1052] <= 12'hfa8; 
COS_ROM[1053] <= 12'hfa5; 
COS_ROM[1054] <= 12'hfa2; 
COS_ROM[1055] <= 12'hf9f; 
COS_ROM[1056] <= 12'hf9c; 
COS_ROM[1057] <= 12'hf98; 
COS_ROM[1058] <= 12'hf95; 
COS_ROM[1059] <= 12'hf92; 
COS_ROM[1060] <= 12'hf8f; 
COS_ROM[1061] <= 12'hf8c; 
COS_ROM[1062] <= 12'hf89; 
COS_ROM[1063] <= 12'hf86; 
COS_ROM[1064] <= 12'hf82; 
COS_ROM[1065] <= 12'hf7f; 
COS_ROM[1066] <= 12'hf7c; 
COS_ROM[1067] <= 12'hf79; 
COS_ROM[1068] <= 12'hf76; 
COS_ROM[1069] <= 12'hf73; 
COS_ROM[1070] <= 12'hf70; 
COS_ROM[1071] <= 12'hf6d; 
COS_ROM[1072] <= 12'hf69; 
COS_ROM[1073] <= 12'hf66; 
COS_ROM[1074] <= 12'hf63; 
COS_ROM[1075] <= 12'hf60; 
COS_ROM[1076] <= 12'hf5d; 
COS_ROM[1077] <= 12'hf5a; 
COS_ROM[1078] <= 12'hf57; 
COS_ROM[1079] <= 12'hf54; 
COS_ROM[1080] <= 12'hf50; 
COS_ROM[1081] <= 12'hf4d; 
COS_ROM[1082] <= 12'hf4a; 
COS_ROM[1083] <= 12'hf47; 
COS_ROM[1084] <= 12'hf44; 
COS_ROM[1085] <= 12'hf41; 
COS_ROM[1086] <= 12'hf3e; 
COS_ROM[1087] <= 12'hf3a; 
COS_ROM[1088] <= 12'hf37; 
COS_ROM[1089] <= 12'hf34; 
COS_ROM[1090] <= 12'hf31; 
COS_ROM[1091] <= 12'hf2e; 
COS_ROM[1092] <= 12'hf2b; 
COS_ROM[1093] <= 12'hf28; 
COS_ROM[1094] <= 12'hf25; 
COS_ROM[1095] <= 12'hf21; 
COS_ROM[1096] <= 12'hf1e; 
COS_ROM[1097] <= 12'hf1b; 
COS_ROM[1098] <= 12'hf18; 
COS_ROM[1099] <= 12'hf15; 
COS_ROM[1100] <= 12'hf12; 
COS_ROM[1101] <= 12'hf0f; 
COS_ROM[1102] <= 12'hf0c; 
COS_ROM[1103] <= 12'hf09; 
COS_ROM[1104] <= 12'hf05; 
COS_ROM[1105] <= 12'hf02; 
COS_ROM[1106] <= 12'heff; 
COS_ROM[1107] <= 12'hefc; 
COS_ROM[1108] <= 12'hef9; 
COS_ROM[1109] <= 12'hef6; 
COS_ROM[1110] <= 12'hef3; 
COS_ROM[1111] <= 12'hef0; 
COS_ROM[1112] <= 12'heed; 
COS_ROM[1113] <= 12'hee9; 
COS_ROM[1114] <= 12'hee6; 
COS_ROM[1115] <= 12'hee3; 
COS_ROM[1116] <= 12'hee0; 
COS_ROM[1117] <= 12'hedd; 
COS_ROM[1118] <= 12'heda; 
COS_ROM[1119] <= 12'hed7; 
COS_ROM[1120] <= 12'hed4; 
COS_ROM[1121] <= 12'hed1; 
COS_ROM[1122] <= 12'hecd; 
COS_ROM[1123] <= 12'heca; 
COS_ROM[1124] <= 12'hec7; 
COS_ROM[1125] <= 12'hec4; 
COS_ROM[1126] <= 12'hec1; 
COS_ROM[1127] <= 12'hebe; 
COS_ROM[1128] <= 12'hebb; 
COS_ROM[1129] <= 12'heb8; 
COS_ROM[1130] <= 12'heb5; 
COS_ROM[1131] <= 12'heb2; 
COS_ROM[1132] <= 12'heae; 
COS_ROM[1133] <= 12'heab; 
COS_ROM[1134] <= 12'hea8; 
COS_ROM[1135] <= 12'hea5; 
COS_ROM[1136] <= 12'hea2; 
COS_ROM[1137] <= 12'he9f; 
COS_ROM[1138] <= 12'he9c; 
COS_ROM[1139] <= 12'he99; 
COS_ROM[1140] <= 12'he96; 
COS_ROM[1141] <= 12'he93; 
COS_ROM[1142] <= 12'he8f; 
COS_ROM[1143] <= 12'he8c; 
COS_ROM[1144] <= 12'he89; 
COS_ROM[1145] <= 12'he86; 
COS_ROM[1146] <= 12'he83; 
COS_ROM[1147] <= 12'he80; 
COS_ROM[1148] <= 12'he7d; 
COS_ROM[1149] <= 12'he7a; 
COS_ROM[1150] <= 12'he77; 
COS_ROM[1151] <= 12'he74; 
COS_ROM[1152] <= 12'he71; 
COS_ROM[1153] <= 12'he6e; 
COS_ROM[1154] <= 12'he6a; 
COS_ROM[1155] <= 12'he67; 
COS_ROM[1156] <= 12'he64; 
COS_ROM[1157] <= 12'he61; 
COS_ROM[1158] <= 12'he5e; 
COS_ROM[1159] <= 12'he5b; 
COS_ROM[1160] <= 12'he58; 
COS_ROM[1161] <= 12'he55; 
COS_ROM[1162] <= 12'he52; 
COS_ROM[1163] <= 12'he4f; 
COS_ROM[1164] <= 12'he4c; 
COS_ROM[1165] <= 12'he49; 
COS_ROM[1166] <= 12'he46; 
COS_ROM[1167] <= 12'he43; 
COS_ROM[1168] <= 12'he3f; 
COS_ROM[1169] <= 12'he3c; 
COS_ROM[1170] <= 12'he39; 
COS_ROM[1171] <= 12'he36; 
COS_ROM[1172] <= 12'he33; 
COS_ROM[1173] <= 12'he30; 
COS_ROM[1174] <= 12'he2d; 
COS_ROM[1175] <= 12'he2a; 
COS_ROM[1176] <= 12'he27; 
COS_ROM[1177] <= 12'he24; 
COS_ROM[1178] <= 12'he21; 
COS_ROM[1179] <= 12'he1e; 
COS_ROM[1180] <= 12'he1b; 
COS_ROM[1181] <= 12'he18; 
COS_ROM[1182] <= 12'he15; 
COS_ROM[1183] <= 12'he12; 
COS_ROM[1184] <= 12'he0f; 
COS_ROM[1185] <= 12'he0c; 
COS_ROM[1186] <= 12'he09; 
COS_ROM[1187] <= 12'he05; 
COS_ROM[1188] <= 12'he02; 
COS_ROM[1189] <= 12'hdff; 
COS_ROM[1190] <= 12'hdfc; 
COS_ROM[1191] <= 12'hdf9; 
COS_ROM[1192] <= 12'hdf6; 
COS_ROM[1193] <= 12'hdf3; 
COS_ROM[1194] <= 12'hdf0; 
COS_ROM[1195] <= 12'hded; 
COS_ROM[1196] <= 12'hdea; 
COS_ROM[1197] <= 12'hde7; 
COS_ROM[1198] <= 12'hde4; 
COS_ROM[1199] <= 12'hde1; 
COS_ROM[1200] <= 12'hdde; 
COS_ROM[1201] <= 12'hddb; 
COS_ROM[1202] <= 12'hdd8; 
COS_ROM[1203] <= 12'hdd5; 
COS_ROM[1204] <= 12'hdd2; 
COS_ROM[1205] <= 12'hdcf; 
COS_ROM[1206] <= 12'hdcc; 
COS_ROM[1207] <= 12'hdc9; 
COS_ROM[1208] <= 12'hdc6; 
COS_ROM[1209] <= 12'hdc3; 
COS_ROM[1210] <= 12'hdc0; 
COS_ROM[1211] <= 12'hdbd; 
COS_ROM[1212] <= 12'hdba; 
COS_ROM[1213] <= 12'hdb7; 
COS_ROM[1214] <= 12'hdb4; 
COS_ROM[1215] <= 12'hdb1; 
COS_ROM[1216] <= 12'hdae; 
COS_ROM[1217] <= 12'hdab; 
COS_ROM[1218] <= 12'hda8; 
COS_ROM[1219] <= 12'hda5; 
COS_ROM[1220] <= 12'hda2; 
COS_ROM[1221] <= 12'hd9f; 
COS_ROM[1222] <= 12'hd9c; 
COS_ROM[1223] <= 12'hd99; 
COS_ROM[1224] <= 12'hd96; 
COS_ROM[1225] <= 12'hd93; 
COS_ROM[1226] <= 12'hd90; 
COS_ROM[1227] <= 12'hd8d; 
COS_ROM[1228] <= 12'hd8a; 
COS_ROM[1229] <= 12'hd87; 
COS_ROM[1230] <= 12'hd84; 
COS_ROM[1231] <= 12'hd81; 
COS_ROM[1232] <= 12'hd7e; 
COS_ROM[1233] <= 12'hd7b; 
COS_ROM[1234] <= 12'hd78; 
COS_ROM[1235] <= 12'hd75; 
COS_ROM[1236] <= 12'hd72; 
COS_ROM[1237] <= 12'hd6f; 
COS_ROM[1238] <= 12'hd6c; 
COS_ROM[1239] <= 12'hd69; 
COS_ROM[1240] <= 12'hd66; 
COS_ROM[1241] <= 12'hd63; 
COS_ROM[1242] <= 12'hd60; 
COS_ROM[1243] <= 12'hd5d; 
COS_ROM[1244] <= 12'hd5a; 
COS_ROM[1245] <= 12'hd57; 
COS_ROM[1246] <= 12'hd54; 
COS_ROM[1247] <= 12'hd51; 
COS_ROM[1248] <= 12'hd4e; 
COS_ROM[1249] <= 12'hd4b; 
COS_ROM[1250] <= 12'hd48; 
COS_ROM[1251] <= 12'hd46; 
COS_ROM[1252] <= 12'hd43; 
COS_ROM[1253] <= 12'hd40; 
COS_ROM[1254] <= 12'hd3d; 
COS_ROM[1255] <= 12'hd3a; 
COS_ROM[1256] <= 12'hd37; 
COS_ROM[1257] <= 12'hd34; 
COS_ROM[1258] <= 12'hd31; 
COS_ROM[1259] <= 12'hd2e; 
COS_ROM[1260] <= 12'hd2b; 
COS_ROM[1261] <= 12'hd28; 
COS_ROM[1262] <= 12'hd25; 
COS_ROM[1263] <= 12'hd22; 
COS_ROM[1264] <= 12'hd1f; 
COS_ROM[1265] <= 12'hd1c; 
COS_ROM[1266] <= 12'hd19; 
COS_ROM[1267] <= 12'hd17; 
COS_ROM[1268] <= 12'hd14; 
COS_ROM[1269] <= 12'hd11; 
COS_ROM[1270] <= 12'hd0e; 
COS_ROM[1271] <= 12'hd0b; 
COS_ROM[1272] <= 12'hd08; 
COS_ROM[1273] <= 12'hd05; 
COS_ROM[1274] <= 12'hd02; 
COS_ROM[1275] <= 12'hcff; 
COS_ROM[1276] <= 12'hcfc; 
COS_ROM[1277] <= 12'hcf9; 
COS_ROM[1278] <= 12'hcf6; 
COS_ROM[1279] <= 12'hcf4; 
COS_ROM[1280] <= 12'hcf1; 
COS_ROM[1281] <= 12'hcee; 
COS_ROM[1282] <= 12'hceb; 
COS_ROM[1283] <= 12'hce8; 
COS_ROM[1284] <= 12'hce5; 
COS_ROM[1285] <= 12'hce2; 
COS_ROM[1286] <= 12'hcdf; 
COS_ROM[1287] <= 12'hcdc; 
COS_ROM[1288] <= 12'hcd9; 
COS_ROM[1289] <= 12'hcd7; 
COS_ROM[1290] <= 12'hcd4; 
COS_ROM[1291] <= 12'hcd1; 
COS_ROM[1292] <= 12'hcce; 
COS_ROM[1293] <= 12'hccb; 
COS_ROM[1294] <= 12'hcc8; 
COS_ROM[1295] <= 12'hcc5; 
COS_ROM[1296] <= 12'hcc2; 
COS_ROM[1297] <= 12'hcc0; 
COS_ROM[1298] <= 12'hcbd; 
COS_ROM[1299] <= 12'hcba; 
COS_ROM[1300] <= 12'hcb7; 
COS_ROM[1301] <= 12'hcb4; 
COS_ROM[1302] <= 12'hcb1; 
COS_ROM[1303] <= 12'hcae; 
COS_ROM[1304] <= 12'hcac; 
COS_ROM[1305] <= 12'hca9; 
COS_ROM[1306] <= 12'hca6; 
COS_ROM[1307] <= 12'hca3; 
COS_ROM[1308] <= 12'hca0; 
COS_ROM[1309] <= 12'hc9d; 
COS_ROM[1310] <= 12'hc9a; 
COS_ROM[1311] <= 12'hc98; 
COS_ROM[1312] <= 12'hc95; 
COS_ROM[1313] <= 12'hc92; 
COS_ROM[1314] <= 12'hc8f; 
COS_ROM[1315] <= 12'hc8c; 
COS_ROM[1316] <= 12'hc89; 
COS_ROM[1317] <= 12'hc87; 
COS_ROM[1318] <= 12'hc84; 
COS_ROM[1319] <= 12'hc81; 
COS_ROM[1320] <= 12'hc7e; 
COS_ROM[1321] <= 12'hc7b; 
COS_ROM[1322] <= 12'hc79; 
COS_ROM[1323] <= 12'hc76; 
COS_ROM[1324] <= 12'hc73; 
COS_ROM[1325] <= 12'hc70; 
COS_ROM[1326] <= 12'hc6d; 
COS_ROM[1327] <= 12'hc6a; 
COS_ROM[1328] <= 12'hc68; 
COS_ROM[1329] <= 12'hc65; 
COS_ROM[1330] <= 12'hc62; 
COS_ROM[1331] <= 12'hc5f; 
COS_ROM[1332] <= 12'hc5c; 
COS_ROM[1333] <= 12'hc5a; 
COS_ROM[1334] <= 12'hc57; 
COS_ROM[1335] <= 12'hc54; 
COS_ROM[1336] <= 12'hc51; 
COS_ROM[1337] <= 12'hc4e; 
COS_ROM[1338] <= 12'hc4c; 
COS_ROM[1339] <= 12'hc49; 
COS_ROM[1340] <= 12'hc46; 
COS_ROM[1341] <= 12'hc43; 
COS_ROM[1342] <= 12'hc41; 
COS_ROM[1343] <= 12'hc3e; 
COS_ROM[1344] <= 12'hc3b; 
COS_ROM[1345] <= 12'hc38; 
COS_ROM[1346] <= 12'hc36; 
COS_ROM[1347] <= 12'hc33; 
COS_ROM[1348] <= 12'hc30; 
COS_ROM[1349] <= 12'hc2d; 
COS_ROM[1350] <= 12'hc2a; 
COS_ROM[1351] <= 12'hc28; 
COS_ROM[1352] <= 12'hc25; 
COS_ROM[1353] <= 12'hc22; 
COS_ROM[1354] <= 12'hc1f; 
COS_ROM[1355] <= 12'hc1d; 
COS_ROM[1356] <= 12'hc1a; 
COS_ROM[1357] <= 12'hc17; 
COS_ROM[1358] <= 12'hc15; 
COS_ROM[1359] <= 12'hc12; 
COS_ROM[1360] <= 12'hc0f; 
COS_ROM[1361] <= 12'hc0c; 
COS_ROM[1362] <= 12'hc0a; 
COS_ROM[1363] <= 12'hc07; 
COS_ROM[1364] <= 12'hc04; 
COS_ROM[1365] <= 12'hc01; 
COS_ROM[1366] <= 12'hbff; 
COS_ROM[1367] <= 12'hbfc; 
COS_ROM[1368] <= 12'hbf9; 
COS_ROM[1369] <= 12'hbf7; 
COS_ROM[1370] <= 12'hbf4; 
COS_ROM[1371] <= 12'hbf1; 
COS_ROM[1372] <= 12'hbee; 
COS_ROM[1373] <= 12'hbec; 
COS_ROM[1374] <= 12'hbe9; 
COS_ROM[1375] <= 12'hbe6; 
COS_ROM[1376] <= 12'hbe4; 
COS_ROM[1377] <= 12'hbe1; 
COS_ROM[1378] <= 12'hbde; 
COS_ROM[1379] <= 12'hbdc; 
COS_ROM[1380] <= 12'hbd9; 
COS_ROM[1381] <= 12'hbd6; 
COS_ROM[1382] <= 12'hbd4; 
COS_ROM[1383] <= 12'hbd1; 
COS_ROM[1384] <= 12'hbce; 
COS_ROM[1385] <= 12'hbcb; 
COS_ROM[1386] <= 12'hbc9; 
COS_ROM[1387] <= 12'hbc6; 
COS_ROM[1388] <= 12'hbc3; 
COS_ROM[1389] <= 12'hbc1; 
COS_ROM[1390] <= 12'hbbe; 
COS_ROM[1391] <= 12'hbbc; 
COS_ROM[1392] <= 12'hbb9; 
COS_ROM[1393] <= 12'hbb6; 
COS_ROM[1394] <= 12'hbb4; 
COS_ROM[1395] <= 12'hbb1; 
COS_ROM[1396] <= 12'hbae; 
COS_ROM[1397] <= 12'hbac; 
COS_ROM[1398] <= 12'hba9; 
COS_ROM[1399] <= 12'hba6; 
COS_ROM[1400] <= 12'hba4; 
COS_ROM[1401] <= 12'hba1; 
COS_ROM[1402] <= 12'hb9e; 
COS_ROM[1403] <= 12'hb9c; 
COS_ROM[1404] <= 12'hb99; 
COS_ROM[1405] <= 12'hb97; 
COS_ROM[1406] <= 12'hb94; 
COS_ROM[1407] <= 12'hb91; 
COS_ROM[1408] <= 12'hb8f; 
COS_ROM[1409] <= 12'hb8c; 
COS_ROM[1410] <= 12'hb8a; 
COS_ROM[1411] <= 12'hb87; 
COS_ROM[1412] <= 12'hb84; 
COS_ROM[1413] <= 12'hb82; 
COS_ROM[1414] <= 12'hb7f; 
COS_ROM[1415] <= 12'hb7d; 
COS_ROM[1416] <= 12'hb7a; 
COS_ROM[1417] <= 12'hb77; 
COS_ROM[1418] <= 12'hb75; 
COS_ROM[1419] <= 12'hb72; 
COS_ROM[1420] <= 12'hb70; 
COS_ROM[1421] <= 12'hb6d; 
COS_ROM[1422] <= 12'hb6a; 
COS_ROM[1423] <= 12'hb68; 
COS_ROM[1424] <= 12'hb65; 
COS_ROM[1425] <= 12'hb63; 
COS_ROM[1426] <= 12'hb60; 
COS_ROM[1427] <= 12'hb5e; 
COS_ROM[1428] <= 12'hb5b; 
COS_ROM[1429] <= 12'hb59; 
COS_ROM[1430] <= 12'hb56; 
COS_ROM[1431] <= 12'hb53; 
COS_ROM[1432] <= 12'hb51; 
COS_ROM[1433] <= 12'hb4e; 
COS_ROM[1434] <= 12'hb4c; 
COS_ROM[1435] <= 12'hb49; 
COS_ROM[1436] <= 12'hb47; 
COS_ROM[1437] <= 12'hb44; 
COS_ROM[1438] <= 12'hb42; 
COS_ROM[1439] <= 12'hb3f; 
COS_ROM[1440] <= 12'hb3d; 
COS_ROM[1441] <= 12'hb3a; 
COS_ROM[1442] <= 12'hb38; 
COS_ROM[1443] <= 12'hb35; 
COS_ROM[1444] <= 12'hb33; 
COS_ROM[1445] <= 12'hb30; 
COS_ROM[1446] <= 12'hb2e; 
COS_ROM[1447] <= 12'hb2b; 
COS_ROM[1448] <= 12'hb29; 
COS_ROM[1449] <= 12'hb26; 
COS_ROM[1450] <= 12'hb24; 
COS_ROM[1451] <= 12'hb21; 
COS_ROM[1452] <= 12'hb1f; 
COS_ROM[1453] <= 12'hb1c; 
COS_ROM[1454] <= 12'hb1a; 
COS_ROM[1455] <= 12'hb17; 
COS_ROM[1456] <= 12'hb15; 
COS_ROM[1457] <= 12'hb12; 
COS_ROM[1458] <= 12'hb10; 
COS_ROM[1459] <= 12'hb0d; 
COS_ROM[1460] <= 12'hb0b; 
COS_ROM[1461] <= 12'hb08; 
COS_ROM[1462] <= 12'hb06; 
COS_ROM[1463] <= 12'hb03; 
COS_ROM[1464] <= 12'hb01; 
COS_ROM[1465] <= 12'hafe; 
COS_ROM[1466] <= 12'hafc; 
COS_ROM[1467] <= 12'hafa; 
COS_ROM[1468] <= 12'haf7; 
COS_ROM[1469] <= 12'haf5; 
COS_ROM[1470] <= 12'haf2; 
COS_ROM[1471] <= 12'haf0; 
COS_ROM[1472] <= 12'haed; 
COS_ROM[1473] <= 12'haeb; 
COS_ROM[1474] <= 12'hae9; 
COS_ROM[1475] <= 12'hae6; 
COS_ROM[1476] <= 12'hae4; 
COS_ROM[1477] <= 12'hae1; 
COS_ROM[1478] <= 12'hadf; 
COS_ROM[1479] <= 12'hadc; 
COS_ROM[1480] <= 12'hada; 
COS_ROM[1481] <= 12'had8; 
COS_ROM[1482] <= 12'had5; 
COS_ROM[1483] <= 12'had3; 
COS_ROM[1484] <= 12'had0; 
COS_ROM[1485] <= 12'hace; 
COS_ROM[1486] <= 12'hacc; 
COS_ROM[1487] <= 12'hac9; 
COS_ROM[1488] <= 12'hac7; 
COS_ROM[1489] <= 12'hac5; 
COS_ROM[1490] <= 12'hac2; 
COS_ROM[1491] <= 12'hac0; 
COS_ROM[1492] <= 12'habd; 
COS_ROM[1493] <= 12'habb; 
COS_ROM[1494] <= 12'hab9; 
COS_ROM[1495] <= 12'hab6; 
COS_ROM[1496] <= 12'hab4; 
COS_ROM[1497] <= 12'hab2; 
COS_ROM[1498] <= 12'haaf; 
COS_ROM[1499] <= 12'haad; 
COS_ROM[1500] <= 12'haab; 
COS_ROM[1501] <= 12'haa8; 
COS_ROM[1502] <= 12'haa6; 
COS_ROM[1503] <= 12'haa4; 
COS_ROM[1504] <= 12'haa1; 
COS_ROM[1505] <= 12'ha9f; 
COS_ROM[1506] <= 12'ha9d; 
COS_ROM[1507] <= 12'ha9a; 
COS_ROM[1508] <= 12'ha98; 
COS_ROM[1509] <= 12'ha96; 
COS_ROM[1510] <= 12'ha93; 
COS_ROM[1511] <= 12'ha91; 
COS_ROM[1512] <= 12'ha8f; 
COS_ROM[1513] <= 12'ha8d; 
COS_ROM[1514] <= 12'ha8a; 
COS_ROM[1515] <= 12'ha88; 
COS_ROM[1516] <= 12'ha86; 
COS_ROM[1517] <= 12'ha83; 
COS_ROM[1518] <= 12'ha81; 
COS_ROM[1519] <= 12'ha7f; 
COS_ROM[1520] <= 12'ha7d; 
COS_ROM[1521] <= 12'ha7a; 
COS_ROM[1522] <= 12'ha78; 
COS_ROM[1523] <= 12'ha76; 
COS_ROM[1524] <= 12'ha73; 
COS_ROM[1525] <= 12'ha71; 
COS_ROM[1526] <= 12'ha6f; 
COS_ROM[1527] <= 12'ha6d; 
COS_ROM[1528] <= 12'ha6a; 
COS_ROM[1529] <= 12'ha68; 
COS_ROM[1530] <= 12'ha66; 
COS_ROM[1531] <= 12'ha64; 
COS_ROM[1532] <= 12'ha61; 
COS_ROM[1533] <= 12'ha5f; 
COS_ROM[1534] <= 12'ha5d; 
COS_ROM[1535] <= 12'ha5b; 
COS_ROM[1536] <= 12'ha59; 
COS_ROM[1537] <= 12'ha56; 
COS_ROM[1538] <= 12'ha54; 
COS_ROM[1539] <= 12'ha52; 
COS_ROM[1540] <= 12'ha50; 
COS_ROM[1541] <= 12'ha4d; 
COS_ROM[1542] <= 12'ha4b; 
COS_ROM[1543] <= 12'ha49; 
COS_ROM[1544] <= 12'ha47; 
COS_ROM[1545] <= 12'ha45; 
COS_ROM[1546] <= 12'ha43; 
COS_ROM[1547] <= 12'ha40; 
COS_ROM[1548] <= 12'ha3e; 
COS_ROM[1549] <= 12'ha3c; 
COS_ROM[1550] <= 12'ha3a; 
COS_ROM[1551] <= 12'ha38; 
COS_ROM[1552] <= 12'ha35; 
COS_ROM[1553] <= 12'ha33; 
COS_ROM[1554] <= 12'ha31; 
COS_ROM[1555] <= 12'ha2f; 
COS_ROM[1556] <= 12'ha2d; 
COS_ROM[1557] <= 12'ha2b; 
COS_ROM[1558] <= 12'ha29; 
COS_ROM[1559] <= 12'ha26; 
COS_ROM[1560] <= 12'ha24; 
COS_ROM[1561] <= 12'ha22; 
COS_ROM[1562] <= 12'ha20; 
COS_ROM[1563] <= 12'ha1e; 
COS_ROM[1564] <= 12'ha1c; 
COS_ROM[1565] <= 12'ha1a; 
COS_ROM[1566] <= 12'ha17; 
COS_ROM[1567] <= 12'ha15; 
COS_ROM[1568] <= 12'ha13; 
COS_ROM[1569] <= 12'ha11; 
COS_ROM[1570] <= 12'ha0f; 
COS_ROM[1571] <= 12'ha0d; 
COS_ROM[1572] <= 12'ha0b; 
COS_ROM[1573] <= 12'ha09; 
COS_ROM[1574] <= 12'ha07; 
COS_ROM[1575] <= 12'ha05; 
COS_ROM[1576] <= 12'ha03; 
COS_ROM[1577] <= 12'ha00; 
COS_ROM[1578] <= 12'h9fe; 
COS_ROM[1579] <= 12'h9fc; 
COS_ROM[1580] <= 12'h9fa; 
COS_ROM[1581] <= 12'h9f8; 
COS_ROM[1582] <= 12'h9f6; 
COS_ROM[1583] <= 12'h9f4; 
COS_ROM[1584] <= 12'h9f2; 
COS_ROM[1585] <= 12'h9f0; 
COS_ROM[1586] <= 12'h9ee; 
COS_ROM[1587] <= 12'h9ec; 
COS_ROM[1588] <= 12'h9ea; 
COS_ROM[1589] <= 12'h9e8; 
COS_ROM[1590] <= 12'h9e6; 
COS_ROM[1591] <= 12'h9e4; 
COS_ROM[1592] <= 12'h9e2; 
COS_ROM[1593] <= 12'h9e0; 
COS_ROM[1594] <= 12'h9de; 
COS_ROM[1595] <= 12'h9dc; 
COS_ROM[1596] <= 12'h9da; 
COS_ROM[1597] <= 12'h9d8; 
COS_ROM[1598] <= 12'h9d6; 
COS_ROM[1599] <= 12'h9d4; 
COS_ROM[1600] <= 12'h9d2; 
COS_ROM[1601] <= 12'h9d0; 
COS_ROM[1602] <= 12'h9ce; 
COS_ROM[1603] <= 12'h9cc; 
COS_ROM[1604] <= 12'h9ca; 
COS_ROM[1605] <= 12'h9c8; 
COS_ROM[1606] <= 12'h9c6; 
COS_ROM[1607] <= 12'h9c4; 
COS_ROM[1608] <= 12'h9c2; 
COS_ROM[1609] <= 12'h9c0; 
COS_ROM[1610] <= 12'h9be; 
COS_ROM[1611] <= 12'h9bc; 
COS_ROM[1612] <= 12'h9ba; 
COS_ROM[1613] <= 12'h9b8; 
COS_ROM[1614] <= 12'h9b6; 
COS_ROM[1615] <= 12'h9b4; 
COS_ROM[1616] <= 12'h9b2; 
COS_ROM[1617] <= 12'h9b0; 
COS_ROM[1618] <= 12'h9ae; 
COS_ROM[1619] <= 12'h9ac; 
COS_ROM[1620] <= 12'h9ab; 
COS_ROM[1621] <= 12'h9a9; 
COS_ROM[1622] <= 12'h9a7; 
COS_ROM[1623] <= 12'h9a5; 
COS_ROM[1624] <= 12'h9a3; 
COS_ROM[1625] <= 12'h9a1; 
COS_ROM[1626] <= 12'h99f; 
COS_ROM[1627] <= 12'h99d; 
COS_ROM[1628] <= 12'h99b; 
COS_ROM[1629] <= 12'h999; 
COS_ROM[1630] <= 12'h998; 
COS_ROM[1631] <= 12'h996; 
COS_ROM[1632] <= 12'h994; 
COS_ROM[1633] <= 12'h992; 
COS_ROM[1634] <= 12'h990; 
COS_ROM[1635] <= 12'h98e; 
COS_ROM[1636] <= 12'h98c; 
COS_ROM[1637] <= 12'h98b; 
COS_ROM[1638] <= 12'h989; 
COS_ROM[1639] <= 12'h987; 
COS_ROM[1640] <= 12'h985; 
COS_ROM[1641] <= 12'h983; 
COS_ROM[1642] <= 12'h981; 
COS_ROM[1643] <= 12'h97f; 
COS_ROM[1644] <= 12'h97e; 
COS_ROM[1645] <= 12'h97c; 
COS_ROM[1646] <= 12'h97a; 
COS_ROM[1647] <= 12'h978; 
COS_ROM[1648] <= 12'h976; 
COS_ROM[1649] <= 12'h975; 
COS_ROM[1650] <= 12'h973; 
COS_ROM[1651] <= 12'h971; 
COS_ROM[1652] <= 12'h96f; 
COS_ROM[1653] <= 12'h96d; 
COS_ROM[1654] <= 12'h96c; 
COS_ROM[1655] <= 12'h96a; 
COS_ROM[1656] <= 12'h968; 
COS_ROM[1657] <= 12'h966; 
COS_ROM[1658] <= 12'h965; 
COS_ROM[1659] <= 12'h963; 
COS_ROM[1660] <= 12'h961; 
COS_ROM[1661] <= 12'h95f; 
COS_ROM[1662] <= 12'h95d; 
COS_ROM[1663] <= 12'h95c; 
COS_ROM[1664] <= 12'h95a; 
COS_ROM[1665] <= 12'h958; 
COS_ROM[1666] <= 12'h957; 
COS_ROM[1667] <= 12'h955; 
COS_ROM[1668] <= 12'h953; 
COS_ROM[1669] <= 12'h951; 
COS_ROM[1670] <= 12'h950; 
COS_ROM[1671] <= 12'h94e; 
COS_ROM[1672] <= 12'h94c; 
COS_ROM[1673] <= 12'h94a; 
COS_ROM[1674] <= 12'h949; 
COS_ROM[1675] <= 12'h947; 
COS_ROM[1676] <= 12'h945; 
COS_ROM[1677] <= 12'h944; 
COS_ROM[1678] <= 12'h942; 
COS_ROM[1679] <= 12'h940; 
COS_ROM[1680] <= 12'h93f; 
COS_ROM[1681] <= 12'h93d; 
COS_ROM[1682] <= 12'h93b; 
COS_ROM[1683] <= 12'h93a; 
COS_ROM[1684] <= 12'h938; 
COS_ROM[1685] <= 12'h936; 
COS_ROM[1686] <= 12'h935; 
COS_ROM[1687] <= 12'h933; 
COS_ROM[1688] <= 12'h931; 
COS_ROM[1689] <= 12'h930; 
COS_ROM[1690] <= 12'h92e; 
COS_ROM[1691] <= 12'h92c; 
COS_ROM[1692] <= 12'h92b; 
COS_ROM[1693] <= 12'h929; 
COS_ROM[1694] <= 12'h927; 
COS_ROM[1695] <= 12'h926; 
COS_ROM[1696] <= 12'h924; 
COS_ROM[1697] <= 12'h923; 
COS_ROM[1698] <= 12'h921; 
COS_ROM[1699] <= 12'h91f; 
COS_ROM[1700] <= 12'h91e; 
COS_ROM[1701] <= 12'h91c; 
COS_ROM[1702] <= 12'h91b; 
COS_ROM[1703] <= 12'h919; 
COS_ROM[1704] <= 12'h917; 
COS_ROM[1705] <= 12'h916; 
COS_ROM[1706] <= 12'h914; 
COS_ROM[1707] <= 12'h913; 
COS_ROM[1708] <= 12'h911; 
COS_ROM[1709] <= 12'h910; 
COS_ROM[1710] <= 12'h90e; 
COS_ROM[1711] <= 12'h90c; 
COS_ROM[1712] <= 12'h90b; 
COS_ROM[1713] <= 12'h909; 
COS_ROM[1714] <= 12'h908; 
COS_ROM[1715] <= 12'h906; 
COS_ROM[1716] <= 12'h905; 
COS_ROM[1717] <= 12'h903; 
COS_ROM[1718] <= 12'h902; 
COS_ROM[1719] <= 12'h900; 
COS_ROM[1720] <= 12'h8ff; 
COS_ROM[1721] <= 12'h8fd; 
COS_ROM[1722] <= 12'h8fc; 
COS_ROM[1723] <= 12'h8fa; 
COS_ROM[1724] <= 12'h8f9; 
COS_ROM[1725] <= 12'h8f7; 
COS_ROM[1726] <= 12'h8f6; 
COS_ROM[1727] <= 12'h8f4; 
COS_ROM[1728] <= 12'h8f3; 
COS_ROM[1729] <= 12'h8f1; 
COS_ROM[1730] <= 12'h8f0; 
COS_ROM[1731] <= 12'h8ee; 
COS_ROM[1732] <= 12'h8ed; 
COS_ROM[1733] <= 12'h8eb; 
COS_ROM[1734] <= 12'h8ea; 
COS_ROM[1735] <= 12'h8e8; 
COS_ROM[1736] <= 12'h8e7; 
COS_ROM[1737] <= 12'h8e6; 
COS_ROM[1738] <= 12'h8e4; 
COS_ROM[1739] <= 12'h8e3; 
COS_ROM[1740] <= 12'h8e1; 
COS_ROM[1741] <= 12'h8e0; 
COS_ROM[1742] <= 12'h8de; 
COS_ROM[1743] <= 12'h8dd; 
COS_ROM[1744] <= 12'h8dc; 
COS_ROM[1745] <= 12'h8da; 
COS_ROM[1746] <= 12'h8d9; 
COS_ROM[1747] <= 12'h8d7; 
COS_ROM[1748] <= 12'h8d6; 
COS_ROM[1749] <= 12'h8d5; 
COS_ROM[1750] <= 12'h8d3; 
COS_ROM[1751] <= 12'h8d2; 
COS_ROM[1752] <= 12'h8d0; 
COS_ROM[1753] <= 12'h8cf; 
COS_ROM[1754] <= 12'h8ce; 
COS_ROM[1755] <= 12'h8cc; 
COS_ROM[1756] <= 12'h8cb; 
COS_ROM[1757] <= 12'h8ca; 
COS_ROM[1758] <= 12'h8c8; 
COS_ROM[1759] <= 12'h8c7; 
COS_ROM[1760] <= 12'h8c6; 
COS_ROM[1761] <= 12'h8c4; 
COS_ROM[1762] <= 12'h8c3; 
COS_ROM[1763] <= 12'h8c2; 
COS_ROM[1764] <= 12'h8c0; 
COS_ROM[1765] <= 12'h8bf; 
COS_ROM[1766] <= 12'h8be; 
COS_ROM[1767] <= 12'h8bc; 
COS_ROM[1768] <= 12'h8bb; 
COS_ROM[1769] <= 12'h8ba; 
COS_ROM[1770] <= 12'h8b8; 
COS_ROM[1771] <= 12'h8b7; 
COS_ROM[1772] <= 12'h8b6; 
COS_ROM[1773] <= 12'h8b4; 
COS_ROM[1774] <= 12'h8b3; 
COS_ROM[1775] <= 12'h8b2; 
COS_ROM[1776] <= 12'h8b1; 
COS_ROM[1777] <= 12'h8af; 
COS_ROM[1778] <= 12'h8ae; 
COS_ROM[1779] <= 12'h8ad; 
COS_ROM[1780] <= 12'h8ac; 
COS_ROM[1781] <= 12'h8aa; 
COS_ROM[1782] <= 12'h8a9; 
COS_ROM[1783] <= 12'h8a8; 
COS_ROM[1784] <= 12'h8a7; 
COS_ROM[1785] <= 12'h8a5; 
COS_ROM[1786] <= 12'h8a4; 
COS_ROM[1787] <= 12'h8a3; 
COS_ROM[1788] <= 12'h8a2; 
COS_ROM[1789] <= 12'h8a0; 
COS_ROM[1790] <= 12'h89f; 
COS_ROM[1791] <= 12'h89e; 
COS_ROM[1792] <= 12'h89d; 
COS_ROM[1793] <= 12'h89c; 
COS_ROM[1794] <= 12'h89a; 
COS_ROM[1795] <= 12'h899; 
COS_ROM[1796] <= 12'h898; 
COS_ROM[1797] <= 12'h897; 
COS_ROM[1798] <= 12'h896; 
COS_ROM[1799] <= 12'h895; 
COS_ROM[1800] <= 12'h893; 
COS_ROM[1801] <= 12'h892; 
COS_ROM[1802] <= 12'h891; 
COS_ROM[1803] <= 12'h890; 
COS_ROM[1804] <= 12'h88f; 
COS_ROM[1805] <= 12'h88e; 
COS_ROM[1806] <= 12'h88c; 
COS_ROM[1807] <= 12'h88b; 
COS_ROM[1808] <= 12'h88a; 
COS_ROM[1809] <= 12'h889; 
COS_ROM[1810] <= 12'h888; 
COS_ROM[1811] <= 12'h887; 
COS_ROM[1812] <= 12'h886; 
COS_ROM[1813] <= 12'h885; 
COS_ROM[1814] <= 12'h883; 
COS_ROM[1815] <= 12'h882; 
COS_ROM[1816] <= 12'h881; 
COS_ROM[1817] <= 12'h880; 
COS_ROM[1818] <= 12'h87f; 
COS_ROM[1819] <= 12'h87e; 
COS_ROM[1820] <= 12'h87d; 
COS_ROM[1821] <= 12'h87c; 
COS_ROM[1822] <= 12'h87b; 
COS_ROM[1823] <= 12'h87a; 
COS_ROM[1824] <= 12'h879; 
COS_ROM[1825] <= 12'h878; 
COS_ROM[1826] <= 12'h877; 
COS_ROM[1827] <= 12'h876; 
COS_ROM[1828] <= 12'h874; 
COS_ROM[1829] <= 12'h873; 
COS_ROM[1830] <= 12'h872; 
COS_ROM[1831] <= 12'h871; 
COS_ROM[1832] <= 12'h870; 
COS_ROM[1833] <= 12'h86f; 
COS_ROM[1834] <= 12'h86e; 
COS_ROM[1835] <= 12'h86d; 
COS_ROM[1836] <= 12'h86c; 
COS_ROM[1837] <= 12'h86b; 
COS_ROM[1838] <= 12'h86a; 
COS_ROM[1839] <= 12'h869; 
COS_ROM[1840] <= 12'h868; 
COS_ROM[1841] <= 12'h867; 
COS_ROM[1842] <= 12'h866; 
COS_ROM[1843] <= 12'h865; 
COS_ROM[1844] <= 12'h864; 
COS_ROM[1845] <= 12'h863; 
COS_ROM[1846] <= 12'h862; 
COS_ROM[1847] <= 12'h862; 
COS_ROM[1848] <= 12'h861; 
COS_ROM[1849] <= 12'h860; 
COS_ROM[1850] <= 12'h85f; 
COS_ROM[1851] <= 12'h85e; 
COS_ROM[1852] <= 12'h85d; 
COS_ROM[1853] <= 12'h85c; 
COS_ROM[1854] <= 12'h85b; 
COS_ROM[1855] <= 12'h85a; 
COS_ROM[1856] <= 12'h859; 
COS_ROM[1857] <= 12'h858; 
COS_ROM[1858] <= 12'h857; 
COS_ROM[1859] <= 12'h856; 
COS_ROM[1860] <= 12'h856; 
COS_ROM[1861] <= 12'h855; 
COS_ROM[1862] <= 12'h854; 
COS_ROM[1863] <= 12'h853; 
COS_ROM[1864] <= 12'h852; 
COS_ROM[1865] <= 12'h851; 
COS_ROM[1866] <= 12'h850; 
COS_ROM[1867] <= 12'h84f; 
COS_ROM[1868] <= 12'h84f; 
COS_ROM[1869] <= 12'h84e; 
COS_ROM[1870] <= 12'h84d; 
COS_ROM[1871] <= 12'h84c; 
COS_ROM[1872] <= 12'h84b; 
COS_ROM[1873] <= 12'h84a; 
COS_ROM[1874] <= 12'h849; 
COS_ROM[1875] <= 12'h849; 
COS_ROM[1876] <= 12'h848; 
COS_ROM[1877] <= 12'h847; 
COS_ROM[1878] <= 12'h846; 
COS_ROM[1879] <= 12'h845; 
COS_ROM[1880] <= 12'h845; 
COS_ROM[1881] <= 12'h844; 
COS_ROM[1882] <= 12'h843; 
COS_ROM[1883] <= 12'h842; 
COS_ROM[1884] <= 12'h841; 
COS_ROM[1885] <= 12'h841; 
COS_ROM[1886] <= 12'h840; 
COS_ROM[1887] <= 12'h83f; 
COS_ROM[1888] <= 12'h83e; 
COS_ROM[1889] <= 12'h83e; 
COS_ROM[1890] <= 12'h83d; 
COS_ROM[1891] <= 12'h83c; 
COS_ROM[1892] <= 12'h83b; 
COS_ROM[1893] <= 12'h83b; 
COS_ROM[1894] <= 12'h83a; 
COS_ROM[1895] <= 12'h839; 
COS_ROM[1896] <= 12'h838; 
COS_ROM[1897] <= 12'h838; 
COS_ROM[1898] <= 12'h837; 
COS_ROM[1899] <= 12'h836; 
COS_ROM[1900] <= 12'h836; 
COS_ROM[1901] <= 12'h835; 
COS_ROM[1902] <= 12'h834; 
COS_ROM[1903] <= 12'h833; 
COS_ROM[1904] <= 12'h833; 
COS_ROM[1905] <= 12'h832; 
COS_ROM[1906] <= 12'h831; 
COS_ROM[1907] <= 12'h831; 
COS_ROM[1908] <= 12'h830; 
COS_ROM[1909] <= 12'h82f; 
COS_ROM[1910] <= 12'h82f; 
COS_ROM[1911] <= 12'h82e; 
COS_ROM[1912] <= 12'h82d; 
COS_ROM[1913] <= 12'h82d; 
COS_ROM[1914] <= 12'h82c; 
COS_ROM[1915] <= 12'h82b; 
COS_ROM[1916] <= 12'h82b; 
COS_ROM[1917] <= 12'h82a; 
COS_ROM[1918] <= 12'h82a; 
COS_ROM[1919] <= 12'h829; 
COS_ROM[1920] <= 12'h828; 
COS_ROM[1921] <= 12'h828; 
COS_ROM[1922] <= 12'h827; 
COS_ROM[1923] <= 12'h827; 
COS_ROM[1924] <= 12'h826; 
COS_ROM[1925] <= 12'h825; 
COS_ROM[1926] <= 12'h825; 
COS_ROM[1927] <= 12'h824; 
COS_ROM[1928] <= 12'h824; 
COS_ROM[1929] <= 12'h823; 
COS_ROM[1930] <= 12'h822; 
COS_ROM[1931] <= 12'h822; 
COS_ROM[1932] <= 12'h821; 
COS_ROM[1933] <= 12'h821; 
COS_ROM[1934] <= 12'h820; 
COS_ROM[1935] <= 12'h820; 
COS_ROM[1936] <= 12'h81f; 
COS_ROM[1937] <= 12'h81f; 
COS_ROM[1938] <= 12'h81e; 
COS_ROM[1939] <= 12'h81e; 
COS_ROM[1940] <= 12'h81d; 
COS_ROM[1941] <= 12'h81d; 
COS_ROM[1942] <= 12'h81c; 
COS_ROM[1943] <= 12'h81b; 
COS_ROM[1944] <= 12'h81b; 
COS_ROM[1945] <= 12'h81a; 
COS_ROM[1946] <= 12'h81a; 
COS_ROM[1947] <= 12'h81a; 
COS_ROM[1948] <= 12'h819; 
COS_ROM[1949] <= 12'h819; 
COS_ROM[1950] <= 12'h818; 
COS_ROM[1951] <= 12'h818; 
COS_ROM[1952] <= 12'h817; 
COS_ROM[1953] <= 12'h817; 
COS_ROM[1954] <= 12'h816; 
COS_ROM[1955] <= 12'h816; 
COS_ROM[1956] <= 12'h815; 
COS_ROM[1957] <= 12'h815; 
COS_ROM[1958] <= 12'h814; 
COS_ROM[1959] <= 12'h814; 
COS_ROM[1960] <= 12'h814; 
COS_ROM[1961] <= 12'h813; 
COS_ROM[1962] <= 12'h813; 
COS_ROM[1963] <= 12'h812; 
COS_ROM[1964] <= 12'h812; 
COS_ROM[1965] <= 12'h812; 
COS_ROM[1966] <= 12'h811; 
COS_ROM[1967] <= 12'h811; 
COS_ROM[1968] <= 12'h810; 
COS_ROM[1969] <= 12'h810; 
COS_ROM[1970] <= 12'h810; 
COS_ROM[1971] <= 12'h80f; 
COS_ROM[1972] <= 12'h80f; 
COS_ROM[1973] <= 12'h80f; 
COS_ROM[1974] <= 12'h80e; 
COS_ROM[1975] <= 12'h80e; 
COS_ROM[1976] <= 12'h80d; 
COS_ROM[1977] <= 12'h80d; 
COS_ROM[1978] <= 12'h80d; 
COS_ROM[1979] <= 12'h80c; 
COS_ROM[1980] <= 12'h80c; 
COS_ROM[1981] <= 12'h80c; 
COS_ROM[1982] <= 12'h80b; 
COS_ROM[1983] <= 12'h80b; 
COS_ROM[1984] <= 12'h80b; 
COS_ROM[1985] <= 12'h80b; 
COS_ROM[1986] <= 12'h80a; 
COS_ROM[1987] <= 12'h80a; 
COS_ROM[1988] <= 12'h80a; 
COS_ROM[1989] <= 12'h809; 
COS_ROM[1990] <= 12'h809; 
COS_ROM[1991] <= 12'h809; 
COS_ROM[1992] <= 12'h809; 
COS_ROM[1993] <= 12'h808; 
COS_ROM[1994] <= 12'h808; 
COS_ROM[1995] <= 12'h808; 
COS_ROM[1996] <= 12'h808; 
COS_ROM[1997] <= 12'h807; 
COS_ROM[1998] <= 12'h807; 
COS_ROM[1999] <= 12'h807; 
COS_ROM[2000] <= 12'h807; 
COS_ROM[2001] <= 12'h806; 
COS_ROM[2002] <= 12'h806; 
COS_ROM[2003] <= 12'h806; 
COS_ROM[2004] <= 12'h806; 
COS_ROM[2005] <= 12'h805; 
COS_ROM[2006] <= 12'h805; 
COS_ROM[2007] <= 12'h805; 
COS_ROM[2008] <= 12'h805; 
COS_ROM[2009] <= 12'h805; 
COS_ROM[2010] <= 12'h804; 
COS_ROM[2011] <= 12'h804; 
COS_ROM[2012] <= 12'h804; 
COS_ROM[2013] <= 12'h804; 
COS_ROM[2014] <= 12'h804; 
COS_ROM[2015] <= 12'h804; 
COS_ROM[2016] <= 12'h803; 
COS_ROM[2017] <= 12'h803; 
COS_ROM[2018] <= 12'h803; 
COS_ROM[2019] <= 12'h803; 
COS_ROM[2020] <= 12'h803; 
COS_ROM[2021] <= 12'h803; 
COS_ROM[2022] <= 12'h803; 
COS_ROM[2023] <= 12'h803; 
COS_ROM[2024] <= 12'h802; 
COS_ROM[2025] <= 12'h802; 
COS_ROM[2026] <= 12'h802; 
COS_ROM[2027] <= 12'h802; 
COS_ROM[2028] <= 12'h802; 
COS_ROM[2029] <= 12'h802; 
COS_ROM[2030] <= 12'h802; 
COS_ROM[2031] <= 12'h802; 
COS_ROM[2032] <= 12'h802; 
COS_ROM[2033] <= 12'h802; 
COS_ROM[2034] <= 12'h801; 
COS_ROM[2035] <= 12'h801; 
COS_ROM[2036] <= 12'h801; 
COS_ROM[2037] <= 12'h801; 
COS_ROM[2038] <= 12'h801; 
COS_ROM[2039] <= 12'h801; 
COS_ROM[2040] <= 12'h801; 
COS_ROM[2041] <= 12'h801; 
COS_ROM[2042] <= 12'h801; 
COS_ROM[2043] <= 12'h801; 
COS_ROM[2044] <= 12'h801; 
COS_ROM[2045] <= 12'h801; 
COS_ROM[2046] <= 12'h801; 
COS_ROM[2047] <= 12'h801; 
COS_ROM[2048] <= 12'h801; 
COS_ROM[2049] <= 12'h801; 
COS_ROM[2050] <= 12'h801; 
COS_ROM[2051] <= 12'h801; 
COS_ROM[2052] <= 12'h801; 
COS_ROM[2053] <= 12'h801; 
COS_ROM[2054] <= 12'h801; 
COS_ROM[2055] <= 12'h801; 
COS_ROM[2056] <= 12'h801; 
COS_ROM[2057] <= 12'h801; 
COS_ROM[2058] <= 12'h801; 
COS_ROM[2059] <= 12'h801; 
COS_ROM[2060] <= 12'h801; 
COS_ROM[2061] <= 12'h801; 
COS_ROM[2062] <= 12'h801; 
COS_ROM[2063] <= 12'h802; 
COS_ROM[2064] <= 12'h802; 
COS_ROM[2065] <= 12'h802; 
COS_ROM[2066] <= 12'h802; 
COS_ROM[2067] <= 12'h802; 
COS_ROM[2068] <= 12'h802; 
COS_ROM[2069] <= 12'h802; 
COS_ROM[2070] <= 12'h802; 
COS_ROM[2071] <= 12'h802; 
COS_ROM[2072] <= 12'h802; 
COS_ROM[2073] <= 12'h803; 
COS_ROM[2074] <= 12'h803; 
COS_ROM[2075] <= 12'h803; 
COS_ROM[2076] <= 12'h803; 
COS_ROM[2077] <= 12'h803; 
COS_ROM[2078] <= 12'h803; 
COS_ROM[2079] <= 12'h803; 
COS_ROM[2080] <= 12'h803; 
COS_ROM[2081] <= 12'h804; 
COS_ROM[2082] <= 12'h804; 
COS_ROM[2083] <= 12'h804; 
COS_ROM[2084] <= 12'h804; 
COS_ROM[2085] <= 12'h804; 
COS_ROM[2086] <= 12'h804; 
COS_ROM[2087] <= 12'h805; 
COS_ROM[2088] <= 12'h805; 
COS_ROM[2089] <= 12'h805; 
COS_ROM[2090] <= 12'h805; 
COS_ROM[2091] <= 12'h805; 
COS_ROM[2092] <= 12'h806; 
COS_ROM[2093] <= 12'h806; 
COS_ROM[2094] <= 12'h806; 
COS_ROM[2095] <= 12'h806; 
COS_ROM[2096] <= 12'h807; 
COS_ROM[2097] <= 12'h807; 
COS_ROM[2098] <= 12'h807; 
COS_ROM[2099] <= 12'h807; 
COS_ROM[2100] <= 12'h808; 
COS_ROM[2101] <= 12'h808; 
COS_ROM[2102] <= 12'h808; 
COS_ROM[2103] <= 12'h808; 
COS_ROM[2104] <= 12'h809; 
COS_ROM[2105] <= 12'h809; 
COS_ROM[2106] <= 12'h809; 
COS_ROM[2107] <= 12'h809; 
COS_ROM[2108] <= 12'h80a; 
COS_ROM[2109] <= 12'h80a; 
COS_ROM[2110] <= 12'h80a; 
COS_ROM[2111] <= 12'h80b; 
COS_ROM[2112] <= 12'h80b; 
COS_ROM[2113] <= 12'h80b; 
COS_ROM[2114] <= 12'h80b; 
COS_ROM[2115] <= 12'h80c; 
COS_ROM[2116] <= 12'h80c; 
COS_ROM[2117] <= 12'h80c; 
COS_ROM[2118] <= 12'h80d; 
COS_ROM[2119] <= 12'h80d; 
COS_ROM[2120] <= 12'h80d; 
COS_ROM[2121] <= 12'h80e; 
COS_ROM[2122] <= 12'h80e; 
COS_ROM[2123] <= 12'h80f; 
COS_ROM[2124] <= 12'h80f; 
COS_ROM[2125] <= 12'h80f; 
COS_ROM[2126] <= 12'h810; 
COS_ROM[2127] <= 12'h810; 
COS_ROM[2128] <= 12'h810; 
COS_ROM[2129] <= 12'h811; 
COS_ROM[2130] <= 12'h811; 
COS_ROM[2131] <= 12'h812; 
COS_ROM[2132] <= 12'h812; 
COS_ROM[2133] <= 12'h812; 
COS_ROM[2134] <= 12'h813; 
COS_ROM[2135] <= 12'h813; 
COS_ROM[2136] <= 12'h814; 
COS_ROM[2137] <= 12'h814; 
COS_ROM[2138] <= 12'h814; 
COS_ROM[2139] <= 12'h815; 
COS_ROM[2140] <= 12'h815; 
COS_ROM[2141] <= 12'h816; 
COS_ROM[2142] <= 12'h816; 
COS_ROM[2143] <= 12'h817; 
COS_ROM[2144] <= 12'h817; 
COS_ROM[2145] <= 12'h818; 
COS_ROM[2146] <= 12'h818; 
COS_ROM[2147] <= 12'h819; 
COS_ROM[2148] <= 12'h819; 
COS_ROM[2149] <= 12'h81a; 
COS_ROM[2150] <= 12'h81a; 
COS_ROM[2151] <= 12'h81a; 
COS_ROM[2152] <= 12'h81b; 
COS_ROM[2153] <= 12'h81b; 
COS_ROM[2154] <= 12'h81c; 
COS_ROM[2155] <= 12'h81d; 
COS_ROM[2156] <= 12'h81d; 
COS_ROM[2157] <= 12'h81e; 
COS_ROM[2158] <= 12'h81e; 
COS_ROM[2159] <= 12'h81f; 
COS_ROM[2160] <= 12'h81f; 
COS_ROM[2161] <= 12'h820; 
COS_ROM[2162] <= 12'h820; 
COS_ROM[2163] <= 12'h821; 
COS_ROM[2164] <= 12'h821; 
COS_ROM[2165] <= 12'h822; 
COS_ROM[2166] <= 12'h822; 
COS_ROM[2167] <= 12'h823; 
COS_ROM[2168] <= 12'h824; 
COS_ROM[2169] <= 12'h824; 
COS_ROM[2170] <= 12'h825; 
COS_ROM[2171] <= 12'h825; 
COS_ROM[2172] <= 12'h826; 
COS_ROM[2173] <= 12'h827; 
COS_ROM[2174] <= 12'h827; 
COS_ROM[2175] <= 12'h828; 
COS_ROM[2176] <= 12'h828; 
COS_ROM[2177] <= 12'h829; 
COS_ROM[2178] <= 12'h82a; 
COS_ROM[2179] <= 12'h82a; 
COS_ROM[2180] <= 12'h82b; 
COS_ROM[2181] <= 12'h82b; 
COS_ROM[2182] <= 12'h82c; 
COS_ROM[2183] <= 12'h82d; 
COS_ROM[2184] <= 12'h82d; 
COS_ROM[2185] <= 12'h82e; 
COS_ROM[2186] <= 12'h82f; 
COS_ROM[2187] <= 12'h82f; 
COS_ROM[2188] <= 12'h830; 
COS_ROM[2189] <= 12'h831; 
COS_ROM[2190] <= 12'h831; 
COS_ROM[2191] <= 12'h832; 
COS_ROM[2192] <= 12'h833; 
COS_ROM[2193] <= 12'h833; 
COS_ROM[2194] <= 12'h834; 
COS_ROM[2195] <= 12'h835; 
COS_ROM[2196] <= 12'h836; 
COS_ROM[2197] <= 12'h836; 
COS_ROM[2198] <= 12'h837; 
COS_ROM[2199] <= 12'h838; 
COS_ROM[2200] <= 12'h838; 
COS_ROM[2201] <= 12'h839; 
COS_ROM[2202] <= 12'h83a; 
COS_ROM[2203] <= 12'h83b; 
COS_ROM[2204] <= 12'h83b; 
COS_ROM[2205] <= 12'h83c; 
COS_ROM[2206] <= 12'h83d; 
COS_ROM[2207] <= 12'h83e; 
COS_ROM[2208] <= 12'h83e; 
COS_ROM[2209] <= 12'h83f; 
COS_ROM[2210] <= 12'h840; 
COS_ROM[2211] <= 12'h841; 
COS_ROM[2212] <= 12'h841; 
COS_ROM[2213] <= 12'h842; 
COS_ROM[2214] <= 12'h843; 
COS_ROM[2215] <= 12'h844; 
COS_ROM[2216] <= 12'h845; 
COS_ROM[2217] <= 12'h845; 
COS_ROM[2218] <= 12'h846; 
COS_ROM[2219] <= 12'h847; 
COS_ROM[2220] <= 12'h848; 
COS_ROM[2221] <= 12'h849; 
COS_ROM[2222] <= 12'h849; 
COS_ROM[2223] <= 12'h84a; 
COS_ROM[2224] <= 12'h84b; 
COS_ROM[2225] <= 12'h84c; 
COS_ROM[2226] <= 12'h84d; 
COS_ROM[2227] <= 12'h84e; 
COS_ROM[2228] <= 12'h84f; 
COS_ROM[2229] <= 12'h84f; 
COS_ROM[2230] <= 12'h850; 
COS_ROM[2231] <= 12'h851; 
COS_ROM[2232] <= 12'h852; 
COS_ROM[2233] <= 12'h853; 
COS_ROM[2234] <= 12'h854; 
COS_ROM[2235] <= 12'h855; 
COS_ROM[2236] <= 12'h856; 
COS_ROM[2237] <= 12'h856; 
COS_ROM[2238] <= 12'h857; 
COS_ROM[2239] <= 12'h858; 
COS_ROM[2240] <= 12'h859; 
COS_ROM[2241] <= 12'h85a; 
COS_ROM[2242] <= 12'h85b; 
COS_ROM[2243] <= 12'h85c; 
COS_ROM[2244] <= 12'h85d; 
COS_ROM[2245] <= 12'h85e; 
COS_ROM[2246] <= 12'h85f; 
COS_ROM[2247] <= 12'h860; 
COS_ROM[2248] <= 12'h861; 
COS_ROM[2249] <= 12'h862; 
COS_ROM[2250] <= 12'h862; 
COS_ROM[2251] <= 12'h863; 
COS_ROM[2252] <= 12'h864; 
COS_ROM[2253] <= 12'h865; 
COS_ROM[2254] <= 12'h866; 
COS_ROM[2255] <= 12'h867; 
COS_ROM[2256] <= 12'h868; 
COS_ROM[2257] <= 12'h869; 
COS_ROM[2258] <= 12'h86a; 
COS_ROM[2259] <= 12'h86b; 
COS_ROM[2260] <= 12'h86c; 
COS_ROM[2261] <= 12'h86d; 
COS_ROM[2262] <= 12'h86e; 
COS_ROM[2263] <= 12'h86f; 
COS_ROM[2264] <= 12'h870; 
COS_ROM[2265] <= 12'h871; 
COS_ROM[2266] <= 12'h872; 
COS_ROM[2267] <= 12'h873; 
COS_ROM[2268] <= 12'h874; 
COS_ROM[2269] <= 12'h876; 
COS_ROM[2270] <= 12'h877; 
COS_ROM[2271] <= 12'h878; 
COS_ROM[2272] <= 12'h879; 
COS_ROM[2273] <= 12'h87a; 
COS_ROM[2274] <= 12'h87b; 
COS_ROM[2275] <= 12'h87c; 
COS_ROM[2276] <= 12'h87d; 
COS_ROM[2277] <= 12'h87e; 
COS_ROM[2278] <= 12'h87f; 
COS_ROM[2279] <= 12'h880; 
COS_ROM[2280] <= 12'h881; 
COS_ROM[2281] <= 12'h882; 
COS_ROM[2282] <= 12'h883; 
COS_ROM[2283] <= 12'h885; 
COS_ROM[2284] <= 12'h886; 
COS_ROM[2285] <= 12'h887; 
COS_ROM[2286] <= 12'h888; 
COS_ROM[2287] <= 12'h889; 
COS_ROM[2288] <= 12'h88a; 
COS_ROM[2289] <= 12'h88b; 
COS_ROM[2290] <= 12'h88c; 
COS_ROM[2291] <= 12'h88e; 
COS_ROM[2292] <= 12'h88f; 
COS_ROM[2293] <= 12'h890; 
COS_ROM[2294] <= 12'h891; 
COS_ROM[2295] <= 12'h892; 
COS_ROM[2296] <= 12'h893; 
COS_ROM[2297] <= 12'h895; 
COS_ROM[2298] <= 12'h896; 
COS_ROM[2299] <= 12'h897; 
COS_ROM[2300] <= 12'h898; 
COS_ROM[2301] <= 12'h899; 
COS_ROM[2302] <= 12'h89a; 
COS_ROM[2303] <= 12'h89c; 
COS_ROM[2304] <= 12'h89d; 
COS_ROM[2305] <= 12'h89e; 
COS_ROM[2306] <= 12'h89f; 
COS_ROM[2307] <= 12'h8a0; 
COS_ROM[2308] <= 12'h8a2; 
COS_ROM[2309] <= 12'h8a3; 
COS_ROM[2310] <= 12'h8a4; 
COS_ROM[2311] <= 12'h8a5; 
COS_ROM[2312] <= 12'h8a7; 
COS_ROM[2313] <= 12'h8a8; 
COS_ROM[2314] <= 12'h8a9; 
COS_ROM[2315] <= 12'h8aa; 
COS_ROM[2316] <= 12'h8ac; 
COS_ROM[2317] <= 12'h8ad; 
COS_ROM[2318] <= 12'h8ae; 
COS_ROM[2319] <= 12'h8af; 
COS_ROM[2320] <= 12'h8b1; 
COS_ROM[2321] <= 12'h8b2; 
COS_ROM[2322] <= 12'h8b3; 
COS_ROM[2323] <= 12'h8b4; 
COS_ROM[2324] <= 12'h8b6; 
COS_ROM[2325] <= 12'h8b7; 
COS_ROM[2326] <= 12'h8b8; 
COS_ROM[2327] <= 12'h8ba; 
COS_ROM[2328] <= 12'h8bb; 
COS_ROM[2329] <= 12'h8bc; 
COS_ROM[2330] <= 12'h8be; 
COS_ROM[2331] <= 12'h8bf; 
COS_ROM[2332] <= 12'h8c0; 
COS_ROM[2333] <= 12'h8c2; 
COS_ROM[2334] <= 12'h8c3; 
COS_ROM[2335] <= 12'h8c4; 
COS_ROM[2336] <= 12'h8c6; 
COS_ROM[2337] <= 12'h8c7; 
COS_ROM[2338] <= 12'h8c8; 
COS_ROM[2339] <= 12'h8ca; 
COS_ROM[2340] <= 12'h8cb; 
COS_ROM[2341] <= 12'h8cc; 
COS_ROM[2342] <= 12'h8ce; 
COS_ROM[2343] <= 12'h8cf; 
COS_ROM[2344] <= 12'h8d0; 
COS_ROM[2345] <= 12'h8d2; 
COS_ROM[2346] <= 12'h8d3; 
COS_ROM[2347] <= 12'h8d5; 
COS_ROM[2348] <= 12'h8d6; 
COS_ROM[2349] <= 12'h8d7; 
COS_ROM[2350] <= 12'h8d9; 
COS_ROM[2351] <= 12'h8da; 
COS_ROM[2352] <= 12'h8dc; 
COS_ROM[2353] <= 12'h8dd; 
COS_ROM[2354] <= 12'h8de; 
COS_ROM[2355] <= 12'h8e0; 
COS_ROM[2356] <= 12'h8e1; 
COS_ROM[2357] <= 12'h8e3; 
COS_ROM[2358] <= 12'h8e4; 
COS_ROM[2359] <= 12'h8e6; 
COS_ROM[2360] <= 12'h8e7; 
COS_ROM[2361] <= 12'h8e8; 
COS_ROM[2362] <= 12'h8ea; 
COS_ROM[2363] <= 12'h8eb; 
COS_ROM[2364] <= 12'h8ed; 
COS_ROM[2365] <= 12'h8ee; 
COS_ROM[2366] <= 12'h8f0; 
COS_ROM[2367] <= 12'h8f1; 
COS_ROM[2368] <= 12'h8f3; 
COS_ROM[2369] <= 12'h8f4; 
COS_ROM[2370] <= 12'h8f6; 
COS_ROM[2371] <= 12'h8f7; 
COS_ROM[2372] <= 12'h8f9; 
COS_ROM[2373] <= 12'h8fa; 
COS_ROM[2374] <= 12'h8fc; 
COS_ROM[2375] <= 12'h8fd; 
COS_ROM[2376] <= 12'h8ff; 
COS_ROM[2377] <= 12'h900; 
COS_ROM[2378] <= 12'h902; 
COS_ROM[2379] <= 12'h903; 
COS_ROM[2380] <= 12'h905; 
COS_ROM[2381] <= 12'h906; 
COS_ROM[2382] <= 12'h908; 
COS_ROM[2383] <= 12'h909; 
COS_ROM[2384] <= 12'h90b; 
COS_ROM[2385] <= 12'h90c; 
COS_ROM[2386] <= 12'h90e; 
COS_ROM[2387] <= 12'h910; 
COS_ROM[2388] <= 12'h911; 
COS_ROM[2389] <= 12'h913; 
COS_ROM[2390] <= 12'h914; 
COS_ROM[2391] <= 12'h916; 
COS_ROM[2392] <= 12'h917; 
COS_ROM[2393] <= 12'h919; 
COS_ROM[2394] <= 12'h91b; 
COS_ROM[2395] <= 12'h91c; 
COS_ROM[2396] <= 12'h91e; 
COS_ROM[2397] <= 12'h91f; 
COS_ROM[2398] <= 12'h921; 
COS_ROM[2399] <= 12'h923; 
COS_ROM[2400] <= 12'h924; 
COS_ROM[2401] <= 12'h926; 
COS_ROM[2402] <= 12'h927; 
COS_ROM[2403] <= 12'h929; 
COS_ROM[2404] <= 12'h92b; 
COS_ROM[2405] <= 12'h92c; 
COS_ROM[2406] <= 12'h92e; 
COS_ROM[2407] <= 12'h930; 
COS_ROM[2408] <= 12'h931; 
COS_ROM[2409] <= 12'h933; 
COS_ROM[2410] <= 12'h935; 
COS_ROM[2411] <= 12'h936; 
COS_ROM[2412] <= 12'h938; 
COS_ROM[2413] <= 12'h93a; 
COS_ROM[2414] <= 12'h93b; 
COS_ROM[2415] <= 12'h93d; 
COS_ROM[2416] <= 12'h93f; 
COS_ROM[2417] <= 12'h940; 
COS_ROM[2418] <= 12'h942; 
COS_ROM[2419] <= 12'h944; 
COS_ROM[2420] <= 12'h945; 
COS_ROM[2421] <= 12'h947; 
COS_ROM[2422] <= 12'h949; 
COS_ROM[2423] <= 12'h94a; 
COS_ROM[2424] <= 12'h94c; 
COS_ROM[2425] <= 12'h94e; 
COS_ROM[2426] <= 12'h950; 
COS_ROM[2427] <= 12'h951; 
COS_ROM[2428] <= 12'h953; 
COS_ROM[2429] <= 12'h955; 
COS_ROM[2430] <= 12'h957; 
COS_ROM[2431] <= 12'h958; 
COS_ROM[2432] <= 12'h95a; 
COS_ROM[2433] <= 12'h95c; 
COS_ROM[2434] <= 12'h95d; 
COS_ROM[2435] <= 12'h95f; 
COS_ROM[2436] <= 12'h961; 
COS_ROM[2437] <= 12'h963; 
COS_ROM[2438] <= 12'h965; 
COS_ROM[2439] <= 12'h966; 
COS_ROM[2440] <= 12'h968; 
COS_ROM[2441] <= 12'h96a; 
COS_ROM[2442] <= 12'h96c; 
COS_ROM[2443] <= 12'h96d; 
COS_ROM[2444] <= 12'h96f; 
COS_ROM[2445] <= 12'h971; 
COS_ROM[2446] <= 12'h973; 
COS_ROM[2447] <= 12'h975; 
COS_ROM[2448] <= 12'h976; 
COS_ROM[2449] <= 12'h978; 
COS_ROM[2450] <= 12'h97a; 
COS_ROM[2451] <= 12'h97c; 
COS_ROM[2452] <= 12'h97e; 
COS_ROM[2453] <= 12'h97f; 
COS_ROM[2454] <= 12'h981; 
COS_ROM[2455] <= 12'h983; 
COS_ROM[2456] <= 12'h985; 
COS_ROM[2457] <= 12'h987; 
COS_ROM[2458] <= 12'h989; 
COS_ROM[2459] <= 12'h98b; 
COS_ROM[2460] <= 12'h98c; 
COS_ROM[2461] <= 12'h98e; 
COS_ROM[2462] <= 12'h990; 
COS_ROM[2463] <= 12'h992; 
COS_ROM[2464] <= 12'h994; 
COS_ROM[2465] <= 12'h996; 
COS_ROM[2466] <= 12'h998; 
COS_ROM[2467] <= 12'h999; 
COS_ROM[2468] <= 12'h99b; 
COS_ROM[2469] <= 12'h99d; 
COS_ROM[2470] <= 12'h99f; 
COS_ROM[2471] <= 12'h9a1; 
COS_ROM[2472] <= 12'h9a3; 
COS_ROM[2473] <= 12'h9a5; 
COS_ROM[2474] <= 12'h9a7; 
COS_ROM[2475] <= 12'h9a9; 
COS_ROM[2476] <= 12'h9ab; 
COS_ROM[2477] <= 12'h9ac; 
COS_ROM[2478] <= 12'h9ae; 
COS_ROM[2479] <= 12'h9b0; 
COS_ROM[2480] <= 12'h9b2; 
COS_ROM[2481] <= 12'h9b4; 
COS_ROM[2482] <= 12'h9b6; 
COS_ROM[2483] <= 12'h9b8; 
COS_ROM[2484] <= 12'h9ba; 
COS_ROM[2485] <= 12'h9bc; 
COS_ROM[2486] <= 12'h9be; 
COS_ROM[2487] <= 12'h9c0; 
COS_ROM[2488] <= 12'h9c2; 
COS_ROM[2489] <= 12'h9c4; 
COS_ROM[2490] <= 12'h9c6; 
COS_ROM[2491] <= 12'h9c8; 
COS_ROM[2492] <= 12'h9ca; 
COS_ROM[2493] <= 12'h9cc; 
COS_ROM[2494] <= 12'h9ce; 
COS_ROM[2495] <= 12'h9d0; 
COS_ROM[2496] <= 12'h9d2; 
COS_ROM[2497] <= 12'h9d4; 
COS_ROM[2498] <= 12'h9d6; 
COS_ROM[2499] <= 12'h9d8; 
COS_ROM[2500] <= 12'h9da; 
COS_ROM[2501] <= 12'h9dc; 
COS_ROM[2502] <= 12'h9de; 
COS_ROM[2503] <= 12'h9e0; 
COS_ROM[2504] <= 12'h9e2; 
COS_ROM[2505] <= 12'h9e4; 
COS_ROM[2506] <= 12'h9e6; 
COS_ROM[2507] <= 12'h9e8; 
COS_ROM[2508] <= 12'h9ea; 
COS_ROM[2509] <= 12'h9ec; 
COS_ROM[2510] <= 12'h9ee; 
COS_ROM[2511] <= 12'h9f0; 
COS_ROM[2512] <= 12'h9f2; 
COS_ROM[2513] <= 12'h9f4; 
COS_ROM[2514] <= 12'h9f6; 
COS_ROM[2515] <= 12'h9f8; 
COS_ROM[2516] <= 12'h9fa; 
COS_ROM[2517] <= 12'h9fc; 
COS_ROM[2518] <= 12'h9fe; 
COS_ROM[2519] <= 12'ha00; 
COS_ROM[2520] <= 12'ha03; 
COS_ROM[2521] <= 12'ha05; 
COS_ROM[2522] <= 12'ha07; 
COS_ROM[2523] <= 12'ha09; 
COS_ROM[2524] <= 12'ha0b; 
COS_ROM[2525] <= 12'ha0d; 
COS_ROM[2526] <= 12'ha0f; 
COS_ROM[2527] <= 12'ha11; 
COS_ROM[2528] <= 12'ha13; 
COS_ROM[2529] <= 12'ha15; 
COS_ROM[2530] <= 12'ha17; 
COS_ROM[2531] <= 12'ha1a; 
COS_ROM[2532] <= 12'ha1c; 
COS_ROM[2533] <= 12'ha1e; 
COS_ROM[2534] <= 12'ha20; 
COS_ROM[2535] <= 12'ha22; 
COS_ROM[2536] <= 12'ha24; 
COS_ROM[2537] <= 12'ha26; 
COS_ROM[2538] <= 12'ha29; 
COS_ROM[2539] <= 12'ha2b; 
COS_ROM[2540] <= 12'ha2d; 
COS_ROM[2541] <= 12'ha2f; 
COS_ROM[2542] <= 12'ha31; 
COS_ROM[2543] <= 12'ha33; 
COS_ROM[2544] <= 12'ha35; 
COS_ROM[2545] <= 12'ha38; 
COS_ROM[2546] <= 12'ha3a; 
COS_ROM[2547] <= 12'ha3c; 
COS_ROM[2548] <= 12'ha3e; 
COS_ROM[2549] <= 12'ha40; 
COS_ROM[2550] <= 12'ha43; 
COS_ROM[2551] <= 12'ha45; 
COS_ROM[2552] <= 12'ha47; 
COS_ROM[2553] <= 12'ha49; 
COS_ROM[2554] <= 12'ha4b; 
COS_ROM[2555] <= 12'ha4d; 
COS_ROM[2556] <= 12'ha50; 
COS_ROM[2557] <= 12'ha52; 
COS_ROM[2558] <= 12'ha54; 
COS_ROM[2559] <= 12'ha56; 
COS_ROM[2560] <= 12'ha59; 
COS_ROM[2561] <= 12'ha5b; 
COS_ROM[2562] <= 12'ha5d; 
COS_ROM[2563] <= 12'ha5f; 
COS_ROM[2564] <= 12'ha61; 
COS_ROM[2565] <= 12'ha64; 
COS_ROM[2566] <= 12'ha66; 
COS_ROM[2567] <= 12'ha68; 
COS_ROM[2568] <= 12'ha6a; 
COS_ROM[2569] <= 12'ha6d; 
COS_ROM[2570] <= 12'ha6f; 
COS_ROM[2571] <= 12'ha71; 
COS_ROM[2572] <= 12'ha73; 
COS_ROM[2573] <= 12'ha76; 
COS_ROM[2574] <= 12'ha78; 
COS_ROM[2575] <= 12'ha7a; 
COS_ROM[2576] <= 12'ha7d; 
COS_ROM[2577] <= 12'ha7f; 
COS_ROM[2578] <= 12'ha81; 
COS_ROM[2579] <= 12'ha83; 
COS_ROM[2580] <= 12'ha86; 
COS_ROM[2581] <= 12'ha88; 
COS_ROM[2582] <= 12'ha8a; 
COS_ROM[2583] <= 12'ha8d; 
COS_ROM[2584] <= 12'ha8f; 
COS_ROM[2585] <= 12'ha91; 
COS_ROM[2586] <= 12'ha93; 
COS_ROM[2587] <= 12'ha96; 
COS_ROM[2588] <= 12'ha98; 
COS_ROM[2589] <= 12'ha9a; 
COS_ROM[2590] <= 12'ha9d; 
COS_ROM[2591] <= 12'ha9f; 
COS_ROM[2592] <= 12'haa1; 
COS_ROM[2593] <= 12'haa4; 
COS_ROM[2594] <= 12'haa6; 
COS_ROM[2595] <= 12'haa8; 
COS_ROM[2596] <= 12'haab; 
COS_ROM[2597] <= 12'haad; 
COS_ROM[2598] <= 12'haaf; 
COS_ROM[2599] <= 12'hab2; 
COS_ROM[2600] <= 12'hab4; 
COS_ROM[2601] <= 12'hab6; 
COS_ROM[2602] <= 12'hab9; 
COS_ROM[2603] <= 12'habb; 
COS_ROM[2604] <= 12'habd; 
COS_ROM[2605] <= 12'hac0; 
COS_ROM[2606] <= 12'hac2; 
COS_ROM[2607] <= 12'hac5; 
COS_ROM[2608] <= 12'hac7; 
COS_ROM[2609] <= 12'hac9; 
COS_ROM[2610] <= 12'hacc; 
COS_ROM[2611] <= 12'hace; 
COS_ROM[2612] <= 12'had0; 
COS_ROM[2613] <= 12'had3; 
COS_ROM[2614] <= 12'had5; 
COS_ROM[2615] <= 12'had8; 
COS_ROM[2616] <= 12'hada; 
COS_ROM[2617] <= 12'hadc; 
COS_ROM[2618] <= 12'hadf; 
COS_ROM[2619] <= 12'hae1; 
COS_ROM[2620] <= 12'hae4; 
COS_ROM[2621] <= 12'hae6; 
COS_ROM[2622] <= 12'hae9; 
COS_ROM[2623] <= 12'haeb; 
COS_ROM[2624] <= 12'haed; 
COS_ROM[2625] <= 12'haf0; 
COS_ROM[2626] <= 12'haf2; 
COS_ROM[2627] <= 12'haf5; 
COS_ROM[2628] <= 12'haf7; 
COS_ROM[2629] <= 12'hafa; 
COS_ROM[2630] <= 12'hafc; 
COS_ROM[2631] <= 12'hafe; 
COS_ROM[2632] <= 12'hb01; 
COS_ROM[2633] <= 12'hb03; 
COS_ROM[2634] <= 12'hb06; 
COS_ROM[2635] <= 12'hb08; 
COS_ROM[2636] <= 12'hb0b; 
COS_ROM[2637] <= 12'hb0d; 
COS_ROM[2638] <= 12'hb10; 
COS_ROM[2639] <= 12'hb12; 
COS_ROM[2640] <= 12'hb15; 
COS_ROM[2641] <= 12'hb17; 
COS_ROM[2642] <= 12'hb1a; 
COS_ROM[2643] <= 12'hb1c; 
COS_ROM[2644] <= 12'hb1f; 
COS_ROM[2645] <= 12'hb21; 
COS_ROM[2646] <= 12'hb24; 
COS_ROM[2647] <= 12'hb26; 
COS_ROM[2648] <= 12'hb29; 
COS_ROM[2649] <= 12'hb2b; 
COS_ROM[2650] <= 12'hb2e; 
COS_ROM[2651] <= 12'hb30; 
COS_ROM[2652] <= 12'hb33; 
COS_ROM[2653] <= 12'hb35; 
COS_ROM[2654] <= 12'hb38; 
COS_ROM[2655] <= 12'hb3a; 
COS_ROM[2656] <= 12'hb3d; 
COS_ROM[2657] <= 12'hb3f; 
COS_ROM[2658] <= 12'hb42; 
COS_ROM[2659] <= 12'hb44; 
COS_ROM[2660] <= 12'hb47; 
COS_ROM[2661] <= 12'hb49; 
COS_ROM[2662] <= 12'hb4c; 
COS_ROM[2663] <= 12'hb4e; 
COS_ROM[2664] <= 12'hb51; 
COS_ROM[2665] <= 12'hb53; 
COS_ROM[2666] <= 12'hb56; 
COS_ROM[2667] <= 12'hb59; 
COS_ROM[2668] <= 12'hb5b; 
COS_ROM[2669] <= 12'hb5e; 
COS_ROM[2670] <= 12'hb60; 
COS_ROM[2671] <= 12'hb63; 
COS_ROM[2672] <= 12'hb65; 
COS_ROM[2673] <= 12'hb68; 
COS_ROM[2674] <= 12'hb6a; 
COS_ROM[2675] <= 12'hb6d; 
COS_ROM[2676] <= 12'hb70; 
COS_ROM[2677] <= 12'hb72; 
COS_ROM[2678] <= 12'hb75; 
COS_ROM[2679] <= 12'hb77; 
COS_ROM[2680] <= 12'hb7a; 
COS_ROM[2681] <= 12'hb7d; 
COS_ROM[2682] <= 12'hb7f; 
COS_ROM[2683] <= 12'hb82; 
COS_ROM[2684] <= 12'hb84; 
COS_ROM[2685] <= 12'hb87; 
COS_ROM[2686] <= 12'hb8a; 
COS_ROM[2687] <= 12'hb8c; 
COS_ROM[2688] <= 12'hb8f; 
COS_ROM[2689] <= 12'hb91; 
COS_ROM[2690] <= 12'hb94; 
COS_ROM[2691] <= 12'hb97; 
COS_ROM[2692] <= 12'hb99; 
COS_ROM[2693] <= 12'hb9c; 
COS_ROM[2694] <= 12'hb9e; 
COS_ROM[2695] <= 12'hba1; 
COS_ROM[2696] <= 12'hba4; 
COS_ROM[2697] <= 12'hba6; 
COS_ROM[2698] <= 12'hba9; 
COS_ROM[2699] <= 12'hbac; 
COS_ROM[2700] <= 12'hbae; 
COS_ROM[2701] <= 12'hbb1; 
COS_ROM[2702] <= 12'hbb4; 
COS_ROM[2703] <= 12'hbb6; 
COS_ROM[2704] <= 12'hbb9; 
COS_ROM[2705] <= 12'hbbc; 
COS_ROM[2706] <= 12'hbbe; 
COS_ROM[2707] <= 12'hbc1; 
COS_ROM[2708] <= 12'hbc3; 
COS_ROM[2709] <= 12'hbc6; 
COS_ROM[2710] <= 12'hbc9; 
COS_ROM[2711] <= 12'hbcb; 
COS_ROM[2712] <= 12'hbce; 
COS_ROM[2713] <= 12'hbd1; 
COS_ROM[2714] <= 12'hbd4; 
COS_ROM[2715] <= 12'hbd6; 
COS_ROM[2716] <= 12'hbd9; 
COS_ROM[2717] <= 12'hbdc; 
COS_ROM[2718] <= 12'hbde; 
COS_ROM[2719] <= 12'hbe1; 
COS_ROM[2720] <= 12'hbe4; 
COS_ROM[2721] <= 12'hbe6; 
COS_ROM[2722] <= 12'hbe9; 
COS_ROM[2723] <= 12'hbec; 
COS_ROM[2724] <= 12'hbee; 
COS_ROM[2725] <= 12'hbf1; 
COS_ROM[2726] <= 12'hbf4; 
COS_ROM[2727] <= 12'hbf7; 
COS_ROM[2728] <= 12'hbf9; 
COS_ROM[2729] <= 12'hbfc; 
COS_ROM[2730] <= 12'hbff; 
COS_ROM[2731] <= 12'hc01; 
COS_ROM[2732] <= 12'hc04; 
COS_ROM[2733] <= 12'hc07; 
COS_ROM[2734] <= 12'hc0a; 
COS_ROM[2735] <= 12'hc0c; 
COS_ROM[2736] <= 12'hc0f; 
COS_ROM[2737] <= 12'hc12; 
COS_ROM[2738] <= 12'hc15; 
COS_ROM[2739] <= 12'hc17; 
COS_ROM[2740] <= 12'hc1a; 
COS_ROM[2741] <= 12'hc1d; 
COS_ROM[2742] <= 12'hc1f; 
COS_ROM[2743] <= 12'hc22; 
COS_ROM[2744] <= 12'hc25; 
COS_ROM[2745] <= 12'hc28; 
COS_ROM[2746] <= 12'hc2a; 
COS_ROM[2747] <= 12'hc2d; 
COS_ROM[2748] <= 12'hc30; 
COS_ROM[2749] <= 12'hc33; 
COS_ROM[2750] <= 12'hc36; 
COS_ROM[2751] <= 12'hc38; 
COS_ROM[2752] <= 12'hc3b; 
COS_ROM[2753] <= 12'hc3e; 
COS_ROM[2754] <= 12'hc41; 
COS_ROM[2755] <= 12'hc43; 
COS_ROM[2756] <= 12'hc46; 
COS_ROM[2757] <= 12'hc49; 
COS_ROM[2758] <= 12'hc4c; 
COS_ROM[2759] <= 12'hc4e; 
COS_ROM[2760] <= 12'hc51; 
COS_ROM[2761] <= 12'hc54; 
COS_ROM[2762] <= 12'hc57; 
COS_ROM[2763] <= 12'hc5a; 
COS_ROM[2764] <= 12'hc5c; 
COS_ROM[2765] <= 12'hc5f; 
COS_ROM[2766] <= 12'hc62; 
COS_ROM[2767] <= 12'hc65; 
COS_ROM[2768] <= 12'hc68; 
COS_ROM[2769] <= 12'hc6a; 
COS_ROM[2770] <= 12'hc6d; 
COS_ROM[2771] <= 12'hc70; 
COS_ROM[2772] <= 12'hc73; 
COS_ROM[2773] <= 12'hc76; 
COS_ROM[2774] <= 12'hc79; 
COS_ROM[2775] <= 12'hc7b; 
COS_ROM[2776] <= 12'hc7e; 
COS_ROM[2777] <= 12'hc81; 
COS_ROM[2778] <= 12'hc84; 
COS_ROM[2779] <= 12'hc87; 
COS_ROM[2780] <= 12'hc89; 
COS_ROM[2781] <= 12'hc8c; 
COS_ROM[2782] <= 12'hc8f; 
COS_ROM[2783] <= 12'hc92; 
COS_ROM[2784] <= 12'hc95; 
COS_ROM[2785] <= 12'hc98; 
COS_ROM[2786] <= 12'hc9a; 
COS_ROM[2787] <= 12'hc9d; 
COS_ROM[2788] <= 12'hca0; 
COS_ROM[2789] <= 12'hca3; 
COS_ROM[2790] <= 12'hca6; 
COS_ROM[2791] <= 12'hca9; 
COS_ROM[2792] <= 12'hcac; 
COS_ROM[2793] <= 12'hcae; 
COS_ROM[2794] <= 12'hcb1; 
COS_ROM[2795] <= 12'hcb4; 
COS_ROM[2796] <= 12'hcb7; 
COS_ROM[2797] <= 12'hcba; 
COS_ROM[2798] <= 12'hcbd; 
COS_ROM[2799] <= 12'hcc0; 
COS_ROM[2800] <= 12'hcc2; 
COS_ROM[2801] <= 12'hcc5; 
COS_ROM[2802] <= 12'hcc8; 
COS_ROM[2803] <= 12'hccb; 
COS_ROM[2804] <= 12'hcce; 
COS_ROM[2805] <= 12'hcd1; 
COS_ROM[2806] <= 12'hcd4; 
COS_ROM[2807] <= 12'hcd7; 
COS_ROM[2808] <= 12'hcd9; 
COS_ROM[2809] <= 12'hcdc; 
COS_ROM[2810] <= 12'hcdf; 
COS_ROM[2811] <= 12'hce2; 
COS_ROM[2812] <= 12'hce5; 
COS_ROM[2813] <= 12'hce8; 
COS_ROM[2814] <= 12'hceb; 
COS_ROM[2815] <= 12'hcee; 
COS_ROM[2816] <= 12'hcf1; 
COS_ROM[2817] <= 12'hcf4; 
COS_ROM[2818] <= 12'hcf6; 
COS_ROM[2819] <= 12'hcf9; 
COS_ROM[2820] <= 12'hcfc; 
COS_ROM[2821] <= 12'hcff; 
COS_ROM[2822] <= 12'hd02; 
COS_ROM[2823] <= 12'hd05; 
COS_ROM[2824] <= 12'hd08; 
COS_ROM[2825] <= 12'hd0b; 
COS_ROM[2826] <= 12'hd0e; 
COS_ROM[2827] <= 12'hd11; 
COS_ROM[2828] <= 12'hd14; 
COS_ROM[2829] <= 12'hd17; 
COS_ROM[2830] <= 12'hd19; 
COS_ROM[2831] <= 12'hd1c; 
COS_ROM[2832] <= 12'hd1f; 
COS_ROM[2833] <= 12'hd22; 
COS_ROM[2834] <= 12'hd25; 
COS_ROM[2835] <= 12'hd28; 
COS_ROM[2836] <= 12'hd2b; 
COS_ROM[2837] <= 12'hd2e; 
COS_ROM[2838] <= 12'hd31; 
COS_ROM[2839] <= 12'hd34; 
COS_ROM[2840] <= 12'hd37; 
COS_ROM[2841] <= 12'hd3a; 
COS_ROM[2842] <= 12'hd3d; 
COS_ROM[2843] <= 12'hd40; 
COS_ROM[2844] <= 12'hd43; 
COS_ROM[2845] <= 12'hd46; 
COS_ROM[2846] <= 12'hd48; 
COS_ROM[2847] <= 12'hd4b; 
COS_ROM[2848] <= 12'hd4e; 
COS_ROM[2849] <= 12'hd51; 
COS_ROM[2850] <= 12'hd54; 
COS_ROM[2851] <= 12'hd57; 
COS_ROM[2852] <= 12'hd5a; 
COS_ROM[2853] <= 12'hd5d; 
COS_ROM[2854] <= 12'hd60; 
COS_ROM[2855] <= 12'hd63; 
COS_ROM[2856] <= 12'hd66; 
COS_ROM[2857] <= 12'hd69; 
COS_ROM[2858] <= 12'hd6c; 
COS_ROM[2859] <= 12'hd6f; 
COS_ROM[2860] <= 12'hd72; 
COS_ROM[2861] <= 12'hd75; 
COS_ROM[2862] <= 12'hd78; 
COS_ROM[2863] <= 12'hd7b; 
COS_ROM[2864] <= 12'hd7e; 
COS_ROM[2865] <= 12'hd81; 
COS_ROM[2866] <= 12'hd84; 
COS_ROM[2867] <= 12'hd87; 
COS_ROM[2868] <= 12'hd8a; 
COS_ROM[2869] <= 12'hd8d; 
COS_ROM[2870] <= 12'hd90; 
COS_ROM[2871] <= 12'hd93; 
COS_ROM[2872] <= 12'hd96; 
COS_ROM[2873] <= 12'hd99; 
COS_ROM[2874] <= 12'hd9c; 
COS_ROM[2875] <= 12'hd9f; 
COS_ROM[2876] <= 12'hda2; 
COS_ROM[2877] <= 12'hda5; 
COS_ROM[2878] <= 12'hda8; 
COS_ROM[2879] <= 12'hdab; 
COS_ROM[2880] <= 12'hdae; 
COS_ROM[2881] <= 12'hdb1; 
COS_ROM[2882] <= 12'hdb4; 
COS_ROM[2883] <= 12'hdb7; 
COS_ROM[2884] <= 12'hdba; 
COS_ROM[2885] <= 12'hdbd; 
COS_ROM[2886] <= 12'hdc0; 
COS_ROM[2887] <= 12'hdc3; 
COS_ROM[2888] <= 12'hdc6; 
COS_ROM[2889] <= 12'hdc9; 
COS_ROM[2890] <= 12'hdcc; 
COS_ROM[2891] <= 12'hdcf; 
COS_ROM[2892] <= 12'hdd2; 
COS_ROM[2893] <= 12'hdd5; 
COS_ROM[2894] <= 12'hdd8; 
COS_ROM[2895] <= 12'hddb; 
COS_ROM[2896] <= 12'hdde; 
COS_ROM[2897] <= 12'hde1; 
COS_ROM[2898] <= 12'hde4; 
COS_ROM[2899] <= 12'hde7; 
COS_ROM[2900] <= 12'hdea; 
COS_ROM[2901] <= 12'hded; 
COS_ROM[2902] <= 12'hdf0; 
COS_ROM[2903] <= 12'hdf3; 
COS_ROM[2904] <= 12'hdf6; 
COS_ROM[2905] <= 12'hdf9; 
COS_ROM[2906] <= 12'hdfc; 
COS_ROM[2907] <= 12'hdff; 
COS_ROM[2908] <= 12'he02; 
COS_ROM[2909] <= 12'he05; 
COS_ROM[2910] <= 12'he09; 
COS_ROM[2911] <= 12'he0c; 
COS_ROM[2912] <= 12'he0f; 
COS_ROM[2913] <= 12'he12; 
COS_ROM[2914] <= 12'he15; 
COS_ROM[2915] <= 12'he18; 
COS_ROM[2916] <= 12'he1b; 
COS_ROM[2917] <= 12'he1e; 
COS_ROM[2918] <= 12'he21; 
COS_ROM[2919] <= 12'he24; 
COS_ROM[2920] <= 12'he27; 
COS_ROM[2921] <= 12'he2a; 
COS_ROM[2922] <= 12'he2d; 
COS_ROM[2923] <= 12'he30; 
COS_ROM[2924] <= 12'he33; 
COS_ROM[2925] <= 12'he36; 
COS_ROM[2926] <= 12'he39; 
COS_ROM[2927] <= 12'he3c; 
COS_ROM[2928] <= 12'he3f; 
COS_ROM[2929] <= 12'he43; 
COS_ROM[2930] <= 12'he46; 
COS_ROM[2931] <= 12'he49; 
COS_ROM[2932] <= 12'he4c; 
COS_ROM[2933] <= 12'he4f; 
COS_ROM[2934] <= 12'he52; 
COS_ROM[2935] <= 12'he55; 
COS_ROM[2936] <= 12'he58; 
COS_ROM[2937] <= 12'he5b; 
COS_ROM[2938] <= 12'he5e; 
COS_ROM[2939] <= 12'he61; 
COS_ROM[2940] <= 12'he64; 
COS_ROM[2941] <= 12'he67; 
COS_ROM[2942] <= 12'he6a; 
COS_ROM[2943] <= 12'he6e; 
COS_ROM[2944] <= 12'he71; 
COS_ROM[2945] <= 12'he74; 
COS_ROM[2946] <= 12'he77; 
COS_ROM[2947] <= 12'he7a; 
COS_ROM[2948] <= 12'he7d; 
COS_ROM[2949] <= 12'he80; 
COS_ROM[2950] <= 12'he83; 
COS_ROM[2951] <= 12'he86; 
COS_ROM[2952] <= 12'he89; 
COS_ROM[2953] <= 12'he8c; 
COS_ROM[2954] <= 12'he8f; 
COS_ROM[2955] <= 12'he93; 
COS_ROM[2956] <= 12'he96; 
COS_ROM[2957] <= 12'he99; 
COS_ROM[2958] <= 12'he9c; 
COS_ROM[2959] <= 12'he9f; 
COS_ROM[2960] <= 12'hea2; 
COS_ROM[2961] <= 12'hea5; 
COS_ROM[2962] <= 12'hea8; 
COS_ROM[2963] <= 12'heab; 
COS_ROM[2964] <= 12'heae; 
COS_ROM[2965] <= 12'heb2; 
COS_ROM[2966] <= 12'heb5; 
COS_ROM[2967] <= 12'heb8; 
COS_ROM[2968] <= 12'hebb; 
COS_ROM[2969] <= 12'hebe; 
COS_ROM[2970] <= 12'hec1; 
COS_ROM[2971] <= 12'hec4; 
COS_ROM[2972] <= 12'hec7; 
COS_ROM[2973] <= 12'heca; 
COS_ROM[2974] <= 12'hecd; 
COS_ROM[2975] <= 12'hed1; 
COS_ROM[2976] <= 12'hed4; 
COS_ROM[2977] <= 12'hed7; 
COS_ROM[2978] <= 12'heda; 
COS_ROM[2979] <= 12'hedd; 
COS_ROM[2980] <= 12'hee0; 
COS_ROM[2981] <= 12'hee3; 
COS_ROM[2982] <= 12'hee6; 
COS_ROM[2983] <= 12'hee9; 
COS_ROM[2984] <= 12'heed; 
COS_ROM[2985] <= 12'hef0; 
COS_ROM[2986] <= 12'hef3; 
COS_ROM[2987] <= 12'hef6; 
COS_ROM[2988] <= 12'hef9; 
COS_ROM[2989] <= 12'hefc; 
COS_ROM[2990] <= 12'heff; 
COS_ROM[2991] <= 12'hf02; 
COS_ROM[2992] <= 12'hf05; 
COS_ROM[2993] <= 12'hf09; 
COS_ROM[2994] <= 12'hf0c; 
COS_ROM[2995] <= 12'hf0f; 
COS_ROM[2996] <= 12'hf12; 
COS_ROM[2997] <= 12'hf15; 
COS_ROM[2998] <= 12'hf18; 
COS_ROM[2999] <= 12'hf1b; 
COS_ROM[3000] <= 12'hf1e; 
COS_ROM[3001] <= 12'hf21; 
COS_ROM[3002] <= 12'hf25; 
COS_ROM[3003] <= 12'hf28; 
COS_ROM[3004] <= 12'hf2b; 
COS_ROM[3005] <= 12'hf2e; 
COS_ROM[3006] <= 12'hf31; 
COS_ROM[3007] <= 12'hf34; 
COS_ROM[3008] <= 12'hf37; 
COS_ROM[3009] <= 12'hf3a; 
COS_ROM[3010] <= 12'hf3e; 
COS_ROM[3011] <= 12'hf41; 
COS_ROM[3012] <= 12'hf44; 
COS_ROM[3013] <= 12'hf47; 
COS_ROM[3014] <= 12'hf4a; 
COS_ROM[3015] <= 12'hf4d; 
COS_ROM[3016] <= 12'hf50; 
COS_ROM[3017] <= 12'hf54; 
COS_ROM[3018] <= 12'hf57; 
COS_ROM[3019] <= 12'hf5a; 
COS_ROM[3020] <= 12'hf5d; 
COS_ROM[3021] <= 12'hf60; 
COS_ROM[3022] <= 12'hf63; 
COS_ROM[3023] <= 12'hf66; 
COS_ROM[3024] <= 12'hf69; 
COS_ROM[3025] <= 12'hf6d; 
COS_ROM[3026] <= 12'hf70; 
COS_ROM[3027] <= 12'hf73; 
COS_ROM[3028] <= 12'hf76; 
COS_ROM[3029] <= 12'hf79; 
COS_ROM[3030] <= 12'hf7c; 
COS_ROM[3031] <= 12'hf7f; 
COS_ROM[3032] <= 12'hf82; 
COS_ROM[3033] <= 12'hf86; 
COS_ROM[3034] <= 12'hf89; 
COS_ROM[3035] <= 12'hf8c; 
COS_ROM[3036] <= 12'hf8f; 
COS_ROM[3037] <= 12'hf92; 
COS_ROM[3038] <= 12'hf95; 
COS_ROM[3039] <= 12'hf98; 
COS_ROM[3040] <= 12'hf9c; 
COS_ROM[3041] <= 12'hf9f; 
COS_ROM[3042] <= 12'hfa2; 
COS_ROM[3043] <= 12'hfa5; 
COS_ROM[3044] <= 12'hfa8; 
COS_ROM[3045] <= 12'hfab; 
COS_ROM[3046] <= 12'hfae; 
COS_ROM[3047] <= 12'hfb2; 
COS_ROM[3048] <= 12'hfb5; 
COS_ROM[3049] <= 12'hfb8; 
COS_ROM[3050] <= 12'hfbb; 
COS_ROM[3051] <= 12'hfbe; 
COS_ROM[3052] <= 12'hfc1; 
COS_ROM[3053] <= 12'hfc4; 
COS_ROM[3054] <= 12'hfc7; 
COS_ROM[3055] <= 12'hfcb; 
COS_ROM[3056] <= 12'hfce; 
COS_ROM[3057] <= 12'hfd1; 
COS_ROM[3058] <= 12'hfd4; 
COS_ROM[3059] <= 12'hfd7; 
COS_ROM[3060] <= 12'hfda; 
COS_ROM[3061] <= 12'hfdd; 
COS_ROM[3062] <= 12'hfe1; 
COS_ROM[3063] <= 12'hfe4; 
COS_ROM[3064] <= 12'hfe7; 
COS_ROM[3065] <= 12'hfea; 
COS_ROM[3066] <= 12'hfed; 
COS_ROM[3067] <= 12'hff0; 
COS_ROM[3068] <= 12'hff3; 
COS_ROM[3069] <= 12'hff7; 
COS_ROM[3070] <= 12'hffa; 
COS_ROM[3071] <= 12'hffd; 
COS_ROM[3072] <= 12'h000; 
COS_ROM[3073] <= 12'h003; 
COS_ROM[3074] <= 12'h006; 
COS_ROM[3075] <= 12'h009; 
COS_ROM[3076] <= 12'h00d; 
COS_ROM[3077] <= 12'h010; 
COS_ROM[3078] <= 12'h013; 
COS_ROM[3079] <= 12'h016; 
COS_ROM[3080] <= 12'h019; 
COS_ROM[3081] <= 12'h01c; 
COS_ROM[3082] <= 12'h01f; 
COS_ROM[3083] <= 12'h023; 
COS_ROM[3084] <= 12'h026; 
COS_ROM[3085] <= 12'h029; 
COS_ROM[3086] <= 12'h02c; 
COS_ROM[3087] <= 12'h02f; 
COS_ROM[3088] <= 12'h032; 
COS_ROM[3089] <= 12'h035; 
COS_ROM[3090] <= 12'h039; 
COS_ROM[3091] <= 12'h03c; 
COS_ROM[3092] <= 12'h03f; 
COS_ROM[3093] <= 12'h042; 
COS_ROM[3094] <= 12'h045; 
COS_ROM[3095] <= 12'h048; 
COS_ROM[3096] <= 12'h04b; 
COS_ROM[3097] <= 12'h04e; 
COS_ROM[3098] <= 12'h052; 
COS_ROM[3099] <= 12'h055; 
COS_ROM[3100] <= 12'h058; 
COS_ROM[3101] <= 12'h05b; 
COS_ROM[3102] <= 12'h05e; 
COS_ROM[3103] <= 12'h061; 
COS_ROM[3104] <= 12'h064; 
COS_ROM[3105] <= 12'h068; 
COS_ROM[3106] <= 12'h06b; 
COS_ROM[3107] <= 12'h06e; 
COS_ROM[3108] <= 12'h071; 
COS_ROM[3109] <= 12'h074; 
COS_ROM[3110] <= 12'h077; 
COS_ROM[3111] <= 12'h07a; 
COS_ROM[3112] <= 12'h07e; 
COS_ROM[3113] <= 12'h081; 
COS_ROM[3114] <= 12'h084; 
COS_ROM[3115] <= 12'h087; 
COS_ROM[3116] <= 12'h08a; 
COS_ROM[3117] <= 12'h08d; 
COS_ROM[3118] <= 12'h090; 
COS_ROM[3119] <= 12'h093; 
COS_ROM[3120] <= 12'h097; 
COS_ROM[3121] <= 12'h09a; 
COS_ROM[3122] <= 12'h09d; 
COS_ROM[3123] <= 12'h0a0; 
COS_ROM[3124] <= 12'h0a3; 
COS_ROM[3125] <= 12'h0a6; 
COS_ROM[3126] <= 12'h0a9; 
COS_ROM[3127] <= 12'h0ac; 
COS_ROM[3128] <= 12'h0b0; 
COS_ROM[3129] <= 12'h0b3; 
COS_ROM[3130] <= 12'h0b6; 
COS_ROM[3131] <= 12'h0b9; 
COS_ROM[3132] <= 12'h0bc; 
COS_ROM[3133] <= 12'h0bf; 
COS_ROM[3134] <= 12'h0c2; 
COS_ROM[3135] <= 12'h0c6; 
COS_ROM[3136] <= 12'h0c9; 
COS_ROM[3137] <= 12'h0cc; 
COS_ROM[3138] <= 12'h0cf; 
COS_ROM[3139] <= 12'h0d2; 
COS_ROM[3140] <= 12'h0d5; 
COS_ROM[3141] <= 12'h0d8; 
COS_ROM[3142] <= 12'h0db; 
COS_ROM[3143] <= 12'h0df; 
COS_ROM[3144] <= 12'h0e2; 
COS_ROM[3145] <= 12'h0e5; 
COS_ROM[3146] <= 12'h0e8; 
COS_ROM[3147] <= 12'h0eb; 
COS_ROM[3148] <= 12'h0ee; 
COS_ROM[3149] <= 12'h0f1; 
COS_ROM[3150] <= 12'h0f4; 
COS_ROM[3151] <= 12'h0f7; 
COS_ROM[3152] <= 12'h0fb; 
COS_ROM[3153] <= 12'h0fe; 
COS_ROM[3154] <= 12'h101; 
COS_ROM[3155] <= 12'h104; 
COS_ROM[3156] <= 12'h107; 
COS_ROM[3157] <= 12'h10a; 
COS_ROM[3158] <= 12'h10d; 
COS_ROM[3159] <= 12'h110; 
COS_ROM[3160] <= 12'h113; 
COS_ROM[3161] <= 12'h117; 
COS_ROM[3162] <= 12'h11a; 
COS_ROM[3163] <= 12'h11d; 
COS_ROM[3164] <= 12'h120; 
COS_ROM[3165] <= 12'h123; 
COS_ROM[3166] <= 12'h126; 
COS_ROM[3167] <= 12'h129; 
COS_ROM[3168] <= 12'h12c; 
COS_ROM[3169] <= 12'h12f; 
COS_ROM[3170] <= 12'h133; 
COS_ROM[3171] <= 12'h136; 
COS_ROM[3172] <= 12'h139; 
COS_ROM[3173] <= 12'h13c; 
COS_ROM[3174] <= 12'h13f; 
COS_ROM[3175] <= 12'h142; 
COS_ROM[3176] <= 12'h145; 
COS_ROM[3177] <= 12'h148; 
COS_ROM[3178] <= 12'h14b; 
COS_ROM[3179] <= 12'h14e; 
COS_ROM[3180] <= 12'h152; 
COS_ROM[3181] <= 12'h155; 
COS_ROM[3182] <= 12'h158; 
COS_ROM[3183] <= 12'h15b; 
COS_ROM[3184] <= 12'h15e; 
COS_ROM[3185] <= 12'h161; 
COS_ROM[3186] <= 12'h164; 
COS_ROM[3187] <= 12'h167; 
COS_ROM[3188] <= 12'h16a; 
COS_ROM[3189] <= 12'h16d; 
COS_ROM[3190] <= 12'h171; 
COS_ROM[3191] <= 12'h174; 
COS_ROM[3192] <= 12'h177; 
COS_ROM[3193] <= 12'h17a; 
COS_ROM[3194] <= 12'h17d; 
COS_ROM[3195] <= 12'h180; 
COS_ROM[3196] <= 12'h183; 
COS_ROM[3197] <= 12'h186; 
COS_ROM[3198] <= 12'h189; 
COS_ROM[3199] <= 12'h18c; 
COS_ROM[3200] <= 12'h18f; 
COS_ROM[3201] <= 12'h192; 
COS_ROM[3202] <= 12'h196; 
COS_ROM[3203] <= 12'h199; 
COS_ROM[3204] <= 12'h19c; 
COS_ROM[3205] <= 12'h19f; 
COS_ROM[3206] <= 12'h1a2; 
COS_ROM[3207] <= 12'h1a5; 
COS_ROM[3208] <= 12'h1a8; 
COS_ROM[3209] <= 12'h1ab; 
COS_ROM[3210] <= 12'h1ae; 
COS_ROM[3211] <= 12'h1b1; 
COS_ROM[3212] <= 12'h1b4; 
COS_ROM[3213] <= 12'h1b7; 
COS_ROM[3214] <= 12'h1ba; 
COS_ROM[3215] <= 12'h1bd; 
COS_ROM[3216] <= 12'h1c1; 
COS_ROM[3217] <= 12'h1c4; 
COS_ROM[3218] <= 12'h1c7; 
COS_ROM[3219] <= 12'h1ca; 
COS_ROM[3220] <= 12'h1cd; 
COS_ROM[3221] <= 12'h1d0; 
COS_ROM[3222] <= 12'h1d3; 
COS_ROM[3223] <= 12'h1d6; 
COS_ROM[3224] <= 12'h1d9; 
COS_ROM[3225] <= 12'h1dc; 
COS_ROM[3226] <= 12'h1df; 
COS_ROM[3227] <= 12'h1e2; 
COS_ROM[3228] <= 12'h1e5; 
COS_ROM[3229] <= 12'h1e8; 
COS_ROM[3230] <= 12'h1eb; 
COS_ROM[3231] <= 12'h1ee; 
COS_ROM[3232] <= 12'h1f1; 
COS_ROM[3233] <= 12'h1f4; 
COS_ROM[3234] <= 12'h1f7; 
COS_ROM[3235] <= 12'h1fb; 
COS_ROM[3236] <= 12'h1fe; 
COS_ROM[3237] <= 12'h201; 
COS_ROM[3238] <= 12'h204; 
COS_ROM[3239] <= 12'h207; 
COS_ROM[3240] <= 12'h20a; 
COS_ROM[3241] <= 12'h20d; 
COS_ROM[3242] <= 12'h210; 
COS_ROM[3243] <= 12'h213; 
COS_ROM[3244] <= 12'h216; 
COS_ROM[3245] <= 12'h219; 
COS_ROM[3246] <= 12'h21c; 
COS_ROM[3247] <= 12'h21f; 
COS_ROM[3248] <= 12'h222; 
COS_ROM[3249] <= 12'h225; 
COS_ROM[3250] <= 12'h228; 
COS_ROM[3251] <= 12'h22b; 
COS_ROM[3252] <= 12'h22e; 
COS_ROM[3253] <= 12'h231; 
COS_ROM[3254] <= 12'h234; 
COS_ROM[3255] <= 12'h237; 
COS_ROM[3256] <= 12'h23a; 
COS_ROM[3257] <= 12'h23d; 
COS_ROM[3258] <= 12'h240; 
COS_ROM[3259] <= 12'h243; 
COS_ROM[3260] <= 12'h246; 
COS_ROM[3261] <= 12'h249; 
COS_ROM[3262] <= 12'h24c; 
COS_ROM[3263] <= 12'h24f; 
COS_ROM[3264] <= 12'h252; 
COS_ROM[3265] <= 12'h255; 
COS_ROM[3266] <= 12'h258; 
COS_ROM[3267] <= 12'h25b; 
COS_ROM[3268] <= 12'h25e; 
COS_ROM[3269] <= 12'h261; 
COS_ROM[3270] <= 12'h264; 
COS_ROM[3271] <= 12'h267; 
COS_ROM[3272] <= 12'h26a; 
COS_ROM[3273] <= 12'h26d; 
COS_ROM[3274] <= 12'h270; 
COS_ROM[3275] <= 12'h273; 
COS_ROM[3276] <= 12'h276; 
COS_ROM[3277] <= 12'h279; 
COS_ROM[3278] <= 12'h27c; 
COS_ROM[3279] <= 12'h27f; 
COS_ROM[3280] <= 12'h282; 
COS_ROM[3281] <= 12'h285; 
COS_ROM[3282] <= 12'h288; 
COS_ROM[3283] <= 12'h28b; 
COS_ROM[3284] <= 12'h28e; 
COS_ROM[3285] <= 12'h291; 
COS_ROM[3286] <= 12'h294; 
COS_ROM[3287] <= 12'h297; 
COS_ROM[3288] <= 12'h29a; 
COS_ROM[3289] <= 12'h29d; 
COS_ROM[3290] <= 12'h2a0; 
COS_ROM[3291] <= 12'h2a3; 
COS_ROM[3292] <= 12'h2a6; 
COS_ROM[3293] <= 12'h2a9; 
COS_ROM[3294] <= 12'h2ac; 
COS_ROM[3295] <= 12'h2af; 
COS_ROM[3296] <= 12'h2b2; 
COS_ROM[3297] <= 12'h2b5; 
COS_ROM[3298] <= 12'h2b8; 
COS_ROM[3299] <= 12'h2ba; 
COS_ROM[3300] <= 12'h2bd; 
COS_ROM[3301] <= 12'h2c0; 
COS_ROM[3302] <= 12'h2c3; 
COS_ROM[3303] <= 12'h2c6; 
COS_ROM[3304] <= 12'h2c9; 
COS_ROM[3305] <= 12'h2cc; 
COS_ROM[3306] <= 12'h2cf; 
COS_ROM[3307] <= 12'h2d2; 
COS_ROM[3308] <= 12'h2d5; 
COS_ROM[3309] <= 12'h2d8; 
COS_ROM[3310] <= 12'h2db; 
COS_ROM[3311] <= 12'h2de; 
COS_ROM[3312] <= 12'h2e1; 
COS_ROM[3313] <= 12'h2e4; 
COS_ROM[3314] <= 12'h2e7; 
COS_ROM[3315] <= 12'h2e9; 
COS_ROM[3316] <= 12'h2ec; 
COS_ROM[3317] <= 12'h2ef; 
COS_ROM[3318] <= 12'h2f2; 
COS_ROM[3319] <= 12'h2f5; 
COS_ROM[3320] <= 12'h2f8; 
COS_ROM[3321] <= 12'h2fb; 
COS_ROM[3322] <= 12'h2fe; 
COS_ROM[3323] <= 12'h301; 
COS_ROM[3324] <= 12'h304; 
COS_ROM[3325] <= 12'h307; 
COS_ROM[3326] <= 12'h30a; 
COS_ROM[3327] <= 12'h30c; 
COS_ROM[3328] <= 12'h30f; 
COS_ROM[3329] <= 12'h312; 
COS_ROM[3330] <= 12'h315; 
COS_ROM[3331] <= 12'h318; 
COS_ROM[3332] <= 12'h31b; 
COS_ROM[3333] <= 12'h31e; 
COS_ROM[3334] <= 12'h321; 
COS_ROM[3335] <= 12'h324; 
COS_ROM[3336] <= 12'h327; 
COS_ROM[3337] <= 12'h329; 
COS_ROM[3338] <= 12'h32c; 
COS_ROM[3339] <= 12'h32f; 
COS_ROM[3340] <= 12'h332; 
COS_ROM[3341] <= 12'h335; 
COS_ROM[3342] <= 12'h338; 
COS_ROM[3343] <= 12'h33b; 
COS_ROM[3344] <= 12'h33e; 
COS_ROM[3345] <= 12'h340; 
COS_ROM[3346] <= 12'h343; 
COS_ROM[3347] <= 12'h346; 
COS_ROM[3348] <= 12'h349; 
COS_ROM[3349] <= 12'h34c; 
COS_ROM[3350] <= 12'h34f; 
COS_ROM[3351] <= 12'h352; 
COS_ROM[3352] <= 12'h354; 
COS_ROM[3353] <= 12'h357; 
COS_ROM[3354] <= 12'h35a; 
COS_ROM[3355] <= 12'h35d; 
COS_ROM[3356] <= 12'h360; 
COS_ROM[3357] <= 12'h363; 
COS_ROM[3358] <= 12'h366; 
COS_ROM[3359] <= 12'h368; 
COS_ROM[3360] <= 12'h36b; 
COS_ROM[3361] <= 12'h36e; 
COS_ROM[3362] <= 12'h371; 
COS_ROM[3363] <= 12'h374; 
COS_ROM[3364] <= 12'h377; 
COS_ROM[3365] <= 12'h379; 
COS_ROM[3366] <= 12'h37c; 
COS_ROM[3367] <= 12'h37f; 
COS_ROM[3368] <= 12'h382; 
COS_ROM[3369] <= 12'h385; 
COS_ROM[3370] <= 12'h387; 
COS_ROM[3371] <= 12'h38a; 
COS_ROM[3372] <= 12'h38d; 
COS_ROM[3373] <= 12'h390; 
COS_ROM[3374] <= 12'h393; 
COS_ROM[3375] <= 12'h396; 
COS_ROM[3376] <= 12'h398; 
COS_ROM[3377] <= 12'h39b; 
COS_ROM[3378] <= 12'h39e; 
COS_ROM[3379] <= 12'h3a1; 
COS_ROM[3380] <= 12'h3a4; 
COS_ROM[3381] <= 12'h3a6; 
COS_ROM[3382] <= 12'h3a9; 
COS_ROM[3383] <= 12'h3ac; 
COS_ROM[3384] <= 12'h3af; 
COS_ROM[3385] <= 12'h3b2; 
COS_ROM[3386] <= 12'h3b4; 
COS_ROM[3387] <= 12'h3b7; 
COS_ROM[3388] <= 12'h3ba; 
COS_ROM[3389] <= 12'h3bd; 
COS_ROM[3390] <= 12'h3bf; 
COS_ROM[3391] <= 12'h3c2; 
COS_ROM[3392] <= 12'h3c5; 
COS_ROM[3393] <= 12'h3c8; 
COS_ROM[3394] <= 12'h3ca; 
COS_ROM[3395] <= 12'h3cd; 
COS_ROM[3396] <= 12'h3d0; 
COS_ROM[3397] <= 12'h3d3; 
COS_ROM[3398] <= 12'h3d6; 
COS_ROM[3399] <= 12'h3d8; 
COS_ROM[3400] <= 12'h3db; 
COS_ROM[3401] <= 12'h3de; 
COS_ROM[3402] <= 12'h3e1; 
COS_ROM[3403] <= 12'h3e3; 
COS_ROM[3404] <= 12'h3e6; 
COS_ROM[3405] <= 12'h3e9; 
COS_ROM[3406] <= 12'h3eb; 
COS_ROM[3407] <= 12'h3ee; 
COS_ROM[3408] <= 12'h3f1; 
COS_ROM[3409] <= 12'h3f4; 
COS_ROM[3410] <= 12'h3f6; 
COS_ROM[3411] <= 12'h3f9; 
COS_ROM[3412] <= 12'h3fc; 
COS_ROM[3413] <= 12'h3ff; 
COS_ROM[3414] <= 12'h401; 
COS_ROM[3415] <= 12'h404; 
COS_ROM[3416] <= 12'h407; 
COS_ROM[3417] <= 12'h409; 
COS_ROM[3418] <= 12'h40c; 
COS_ROM[3419] <= 12'h40f; 
COS_ROM[3420] <= 12'h412; 
COS_ROM[3421] <= 12'h414; 
COS_ROM[3422] <= 12'h417; 
COS_ROM[3423] <= 12'h41a; 
COS_ROM[3424] <= 12'h41c; 
COS_ROM[3425] <= 12'h41f; 
COS_ROM[3426] <= 12'h422; 
COS_ROM[3427] <= 12'h424; 
COS_ROM[3428] <= 12'h427; 
COS_ROM[3429] <= 12'h42a; 
COS_ROM[3430] <= 12'h42c; 
COS_ROM[3431] <= 12'h42f; 
COS_ROM[3432] <= 12'h432; 
COS_ROM[3433] <= 12'h435; 
COS_ROM[3434] <= 12'h437; 
COS_ROM[3435] <= 12'h43a; 
COS_ROM[3436] <= 12'h43d; 
COS_ROM[3437] <= 12'h43f; 
COS_ROM[3438] <= 12'h442; 
COS_ROM[3439] <= 12'h444; 
COS_ROM[3440] <= 12'h447; 
COS_ROM[3441] <= 12'h44a; 
COS_ROM[3442] <= 12'h44c; 
COS_ROM[3443] <= 12'h44f; 
COS_ROM[3444] <= 12'h452; 
COS_ROM[3445] <= 12'h454; 
COS_ROM[3446] <= 12'h457; 
COS_ROM[3447] <= 12'h45a; 
COS_ROM[3448] <= 12'h45c; 
COS_ROM[3449] <= 12'h45f; 
COS_ROM[3450] <= 12'h462; 
COS_ROM[3451] <= 12'h464; 
COS_ROM[3452] <= 12'h467; 
COS_ROM[3453] <= 12'h469; 
COS_ROM[3454] <= 12'h46c; 
COS_ROM[3455] <= 12'h46f; 
COS_ROM[3456] <= 12'h471; 
COS_ROM[3457] <= 12'h474; 
COS_ROM[3458] <= 12'h476; 
COS_ROM[3459] <= 12'h479; 
COS_ROM[3460] <= 12'h47c; 
COS_ROM[3461] <= 12'h47e; 
COS_ROM[3462] <= 12'h481; 
COS_ROM[3463] <= 12'h483; 
COS_ROM[3464] <= 12'h486; 
COS_ROM[3465] <= 12'h489; 
COS_ROM[3466] <= 12'h48b; 
COS_ROM[3467] <= 12'h48e; 
COS_ROM[3468] <= 12'h490; 
COS_ROM[3469] <= 12'h493; 
COS_ROM[3470] <= 12'h496; 
COS_ROM[3471] <= 12'h498; 
COS_ROM[3472] <= 12'h49b; 
COS_ROM[3473] <= 12'h49d; 
COS_ROM[3474] <= 12'h4a0; 
COS_ROM[3475] <= 12'h4a2; 
COS_ROM[3476] <= 12'h4a5; 
COS_ROM[3477] <= 12'h4a7; 
COS_ROM[3478] <= 12'h4aa; 
COS_ROM[3479] <= 12'h4ad; 
COS_ROM[3480] <= 12'h4af; 
COS_ROM[3481] <= 12'h4b2; 
COS_ROM[3482] <= 12'h4b4; 
COS_ROM[3483] <= 12'h4b7; 
COS_ROM[3484] <= 12'h4b9; 
COS_ROM[3485] <= 12'h4bc; 
COS_ROM[3486] <= 12'h4be; 
COS_ROM[3487] <= 12'h4c1; 
COS_ROM[3488] <= 12'h4c3; 
COS_ROM[3489] <= 12'h4c6; 
COS_ROM[3490] <= 12'h4c8; 
COS_ROM[3491] <= 12'h4cb; 
COS_ROM[3492] <= 12'h4cd; 
COS_ROM[3493] <= 12'h4d0; 
COS_ROM[3494] <= 12'h4d2; 
COS_ROM[3495] <= 12'h4d5; 
COS_ROM[3496] <= 12'h4d7; 
COS_ROM[3497] <= 12'h4da; 
COS_ROM[3498] <= 12'h4dc; 
COS_ROM[3499] <= 12'h4df; 
COS_ROM[3500] <= 12'h4e1; 
COS_ROM[3501] <= 12'h4e4; 
COS_ROM[3502] <= 12'h4e6; 
COS_ROM[3503] <= 12'h4e9; 
COS_ROM[3504] <= 12'h4eb; 
COS_ROM[3505] <= 12'h4ee; 
COS_ROM[3506] <= 12'h4f0; 
COS_ROM[3507] <= 12'h4f3; 
COS_ROM[3508] <= 12'h4f5; 
COS_ROM[3509] <= 12'h4f8; 
COS_ROM[3510] <= 12'h4fa; 
COS_ROM[3511] <= 12'h4fd; 
COS_ROM[3512] <= 12'h4ff; 
COS_ROM[3513] <= 12'h502; 
COS_ROM[3514] <= 12'h504; 
COS_ROM[3515] <= 12'h506; 
COS_ROM[3516] <= 12'h509; 
COS_ROM[3517] <= 12'h50b; 
COS_ROM[3518] <= 12'h50e; 
COS_ROM[3519] <= 12'h510; 
COS_ROM[3520] <= 12'h513; 
COS_ROM[3521] <= 12'h515; 
COS_ROM[3522] <= 12'h517; 
COS_ROM[3523] <= 12'h51a; 
COS_ROM[3524] <= 12'h51c; 
COS_ROM[3525] <= 12'h51f; 
COS_ROM[3526] <= 12'h521; 
COS_ROM[3527] <= 12'h524; 
COS_ROM[3528] <= 12'h526; 
COS_ROM[3529] <= 12'h528; 
COS_ROM[3530] <= 12'h52b; 
COS_ROM[3531] <= 12'h52d; 
COS_ROM[3532] <= 12'h530; 
COS_ROM[3533] <= 12'h532; 
COS_ROM[3534] <= 12'h534; 
COS_ROM[3535] <= 12'h537; 
COS_ROM[3536] <= 12'h539; 
COS_ROM[3537] <= 12'h53b; 
COS_ROM[3538] <= 12'h53e; 
COS_ROM[3539] <= 12'h540; 
COS_ROM[3540] <= 12'h543; 
COS_ROM[3541] <= 12'h545; 
COS_ROM[3542] <= 12'h547; 
COS_ROM[3543] <= 12'h54a; 
COS_ROM[3544] <= 12'h54c; 
COS_ROM[3545] <= 12'h54e; 
COS_ROM[3546] <= 12'h551; 
COS_ROM[3547] <= 12'h553; 
COS_ROM[3548] <= 12'h555; 
COS_ROM[3549] <= 12'h558; 
COS_ROM[3550] <= 12'h55a; 
COS_ROM[3551] <= 12'h55c; 
COS_ROM[3552] <= 12'h55f; 
COS_ROM[3553] <= 12'h561; 
COS_ROM[3554] <= 12'h563; 
COS_ROM[3555] <= 12'h566; 
COS_ROM[3556] <= 12'h568; 
COS_ROM[3557] <= 12'h56a; 
COS_ROM[3558] <= 12'h56d; 
COS_ROM[3559] <= 12'h56f; 
COS_ROM[3560] <= 12'h571; 
COS_ROM[3561] <= 12'h573; 
COS_ROM[3562] <= 12'h576; 
COS_ROM[3563] <= 12'h578; 
COS_ROM[3564] <= 12'h57a; 
COS_ROM[3565] <= 12'h57d; 
COS_ROM[3566] <= 12'h57f; 
COS_ROM[3567] <= 12'h581; 
COS_ROM[3568] <= 12'h583; 
COS_ROM[3569] <= 12'h586; 
COS_ROM[3570] <= 12'h588; 
COS_ROM[3571] <= 12'h58a; 
COS_ROM[3572] <= 12'h58d; 
COS_ROM[3573] <= 12'h58f; 
COS_ROM[3574] <= 12'h591; 
COS_ROM[3575] <= 12'h593; 
COS_ROM[3576] <= 12'h596; 
COS_ROM[3577] <= 12'h598; 
COS_ROM[3578] <= 12'h59a; 
COS_ROM[3579] <= 12'h59c; 
COS_ROM[3580] <= 12'h59f; 
COS_ROM[3581] <= 12'h5a1; 
COS_ROM[3582] <= 12'h5a3; 
COS_ROM[3583] <= 12'h5a5; 
COS_ROM[3584] <= 12'h5a7; 
COS_ROM[3585] <= 12'h5aa; 
COS_ROM[3586] <= 12'h5ac; 
COS_ROM[3587] <= 12'h5ae; 
COS_ROM[3588] <= 12'h5b0; 
COS_ROM[3589] <= 12'h5b3; 
COS_ROM[3590] <= 12'h5b5; 
COS_ROM[3591] <= 12'h5b7; 
COS_ROM[3592] <= 12'h5b9; 
COS_ROM[3593] <= 12'h5bb; 
COS_ROM[3594] <= 12'h5bd; 
COS_ROM[3595] <= 12'h5c0; 
COS_ROM[3596] <= 12'h5c2; 
COS_ROM[3597] <= 12'h5c4; 
COS_ROM[3598] <= 12'h5c6; 
COS_ROM[3599] <= 12'h5c8; 
COS_ROM[3600] <= 12'h5cb; 
COS_ROM[3601] <= 12'h5cd; 
COS_ROM[3602] <= 12'h5cf; 
COS_ROM[3603] <= 12'h5d1; 
COS_ROM[3604] <= 12'h5d3; 
COS_ROM[3605] <= 12'h5d5; 
COS_ROM[3606] <= 12'h5d7; 
COS_ROM[3607] <= 12'h5da; 
COS_ROM[3608] <= 12'h5dc; 
COS_ROM[3609] <= 12'h5de; 
COS_ROM[3610] <= 12'h5e0; 
COS_ROM[3611] <= 12'h5e2; 
COS_ROM[3612] <= 12'h5e4; 
COS_ROM[3613] <= 12'h5e6; 
COS_ROM[3614] <= 12'h5e9; 
COS_ROM[3615] <= 12'h5eb; 
COS_ROM[3616] <= 12'h5ed; 
COS_ROM[3617] <= 12'h5ef; 
COS_ROM[3618] <= 12'h5f1; 
COS_ROM[3619] <= 12'h5f3; 
COS_ROM[3620] <= 12'h5f5; 
COS_ROM[3621] <= 12'h5f7; 
COS_ROM[3622] <= 12'h5f9; 
COS_ROM[3623] <= 12'h5fb; 
COS_ROM[3624] <= 12'h5fd; 
COS_ROM[3625] <= 12'h600; 
COS_ROM[3626] <= 12'h602; 
COS_ROM[3627] <= 12'h604; 
COS_ROM[3628] <= 12'h606; 
COS_ROM[3629] <= 12'h608; 
COS_ROM[3630] <= 12'h60a; 
COS_ROM[3631] <= 12'h60c; 
COS_ROM[3632] <= 12'h60e; 
COS_ROM[3633] <= 12'h610; 
COS_ROM[3634] <= 12'h612; 
COS_ROM[3635] <= 12'h614; 
COS_ROM[3636] <= 12'h616; 
COS_ROM[3637] <= 12'h618; 
COS_ROM[3638] <= 12'h61a; 
COS_ROM[3639] <= 12'h61c; 
COS_ROM[3640] <= 12'h61e; 
COS_ROM[3641] <= 12'h620; 
COS_ROM[3642] <= 12'h622; 
COS_ROM[3643] <= 12'h624; 
COS_ROM[3644] <= 12'h626; 
COS_ROM[3645] <= 12'h628; 
COS_ROM[3646] <= 12'h62a; 
COS_ROM[3647] <= 12'h62c; 
COS_ROM[3648] <= 12'h62e; 
COS_ROM[3649] <= 12'h630; 
COS_ROM[3650] <= 12'h632; 
COS_ROM[3651] <= 12'h634; 
COS_ROM[3652] <= 12'h636; 
COS_ROM[3653] <= 12'h638; 
COS_ROM[3654] <= 12'h63a; 
COS_ROM[3655] <= 12'h63c; 
COS_ROM[3656] <= 12'h63e; 
COS_ROM[3657] <= 12'h640; 
COS_ROM[3658] <= 12'h642; 
COS_ROM[3659] <= 12'h644; 
COS_ROM[3660] <= 12'h646; 
COS_ROM[3661] <= 12'h648; 
COS_ROM[3662] <= 12'h64a; 
COS_ROM[3663] <= 12'h64c; 
COS_ROM[3664] <= 12'h64e; 
COS_ROM[3665] <= 12'h650; 
COS_ROM[3666] <= 12'h652; 
COS_ROM[3667] <= 12'h654; 
COS_ROM[3668] <= 12'h655; 
COS_ROM[3669] <= 12'h657; 
COS_ROM[3670] <= 12'h659; 
COS_ROM[3671] <= 12'h65b; 
COS_ROM[3672] <= 12'h65d; 
COS_ROM[3673] <= 12'h65f; 
COS_ROM[3674] <= 12'h661; 
COS_ROM[3675] <= 12'h663; 
COS_ROM[3676] <= 12'h665; 
COS_ROM[3677] <= 12'h667; 
COS_ROM[3678] <= 12'h668; 
COS_ROM[3679] <= 12'h66a; 
COS_ROM[3680] <= 12'h66c; 
COS_ROM[3681] <= 12'h66e; 
COS_ROM[3682] <= 12'h670; 
COS_ROM[3683] <= 12'h672; 
COS_ROM[3684] <= 12'h674; 
COS_ROM[3685] <= 12'h675; 
COS_ROM[3686] <= 12'h677; 
COS_ROM[3687] <= 12'h679; 
COS_ROM[3688] <= 12'h67b; 
COS_ROM[3689] <= 12'h67d; 
COS_ROM[3690] <= 12'h67f; 
COS_ROM[3691] <= 12'h681; 
COS_ROM[3692] <= 12'h682; 
COS_ROM[3693] <= 12'h684; 
COS_ROM[3694] <= 12'h686; 
COS_ROM[3695] <= 12'h688; 
COS_ROM[3696] <= 12'h68a; 
COS_ROM[3697] <= 12'h68b; 
COS_ROM[3698] <= 12'h68d; 
COS_ROM[3699] <= 12'h68f; 
COS_ROM[3700] <= 12'h691; 
COS_ROM[3701] <= 12'h693; 
COS_ROM[3702] <= 12'h694; 
COS_ROM[3703] <= 12'h696; 
COS_ROM[3704] <= 12'h698; 
COS_ROM[3705] <= 12'h69a; 
COS_ROM[3706] <= 12'h69b; 
COS_ROM[3707] <= 12'h69d; 
COS_ROM[3708] <= 12'h69f; 
COS_ROM[3709] <= 12'h6a1; 
COS_ROM[3710] <= 12'h6a3; 
COS_ROM[3711] <= 12'h6a4; 
COS_ROM[3712] <= 12'h6a6; 
COS_ROM[3713] <= 12'h6a8; 
COS_ROM[3714] <= 12'h6a9; 
COS_ROM[3715] <= 12'h6ab; 
COS_ROM[3716] <= 12'h6ad; 
COS_ROM[3717] <= 12'h6af; 
COS_ROM[3718] <= 12'h6b0; 
COS_ROM[3719] <= 12'h6b2; 
COS_ROM[3720] <= 12'h6b4; 
COS_ROM[3721] <= 12'h6b6; 
COS_ROM[3722] <= 12'h6b7; 
COS_ROM[3723] <= 12'h6b9; 
COS_ROM[3724] <= 12'h6bb; 
COS_ROM[3725] <= 12'h6bc; 
COS_ROM[3726] <= 12'h6be; 
COS_ROM[3727] <= 12'h6c0; 
COS_ROM[3728] <= 12'h6c1; 
COS_ROM[3729] <= 12'h6c3; 
COS_ROM[3730] <= 12'h6c5; 
COS_ROM[3731] <= 12'h6c6; 
COS_ROM[3732] <= 12'h6c8; 
COS_ROM[3733] <= 12'h6ca; 
COS_ROM[3734] <= 12'h6cb; 
COS_ROM[3735] <= 12'h6cd; 
COS_ROM[3736] <= 12'h6cf; 
COS_ROM[3737] <= 12'h6d0; 
COS_ROM[3738] <= 12'h6d2; 
COS_ROM[3739] <= 12'h6d4; 
COS_ROM[3740] <= 12'h6d5; 
COS_ROM[3741] <= 12'h6d7; 
COS_ROM[3742] <= 12'h6d9; 
COS_ROM[3743] <= 12'h6da; 
COS_ROM[3744] <= 12'h6dc; 
COS_ROM[3745] <= 12'h6dd; 
COS_ROM[3746] <= 12'h6df; 
COS_ROM[3747] <= 12'h6e1; 
COS_ROM[3748] <= 12'h6e2; 
COS_ROM[3749] <= 12'h6e4; 
COS_ROM[3750] <= 12'h6e5; 
COS_ROM[3751] <= 12'h6e7; 
COS_ROM[3752] <= 12'h6e9; 
COS_ROM[3753] <= 12'h6ea; 
COS_ROM[3754] <= 12'h6ec; 
COS_ROM[3755] <= 12'h6ed; 
COS_ROM[3756] <= 12'h6ef; 
COS_ROM[3757] <= 12'h6f0; 
COS_ROM[3758] <= 12'h6f2; 
COS_ROM[3759] <= 12'h6f4; 
COS_ROM[3760] <= 12'h6f5; 
COS_ROM[3761] <= 12'h6f7; 
COS_ROM[3762] <= 12'h6f8; 
COS_ROM[3763] <= 12'h6fa; 
COS_ROM[3764] <= 12'h6fb; 
COS_ROM[3765] <= 12'h6fd; 
COS_ROM[3766] <= 12'h6fe; 
COS_ROM[3767] <= 12'h700; 
COS_ROM[3768] <= 12'h701; 
COS_ROM[3769] <= 12'h703; 
COS_ROM[3770] <= 12'h704; 
COS_ROM[3771] <= 12'h706; 
COS_ROM[3772] <= 12'h707; 
COS_ROM[3773] <= 12'h709; 
COS_ROM[3774] <= 12'h70a; 
COS_ROM[3775] <= 12'h70c; 
COS_ROM[3776] <= 12'h70d; 
COS_ROM[3777] <= 12'h70f; 
COS_ROM[3778] <= 12'h710; 
COS_ROM[3779] <= 12'h712; 
COS_ROM[3780] <= 12'h713; 
COS_ROM[3781] <= 12'h715; 
COS_ROM[3782] <= 12'h716; 
COS_ROM[3783] <= 12'h718; 
COS_ROM[3784] <= 12'h719; 
COS_ROM[3785] <= 12'h71a; 
COS_ROM[3786] <= 12'h71c; 
COS_ROM[3787] <= 12'h71d; 
COS_ROM[3788] <= 12'h71f; 
COS_ROM[3789] <= 12'h720; 
COS_ROM[3790] <= 12'h722; 
COS_ROM[3791] <= 12'h723; 
COS_ROM[3792] <= 12'h724; 
COS_ROM[3793] <= 12'h726; 
COS_ROM[3794] <= 12'h727; 
COS_ROM[3795] <= 12'h729; 
COS_ROM[3796] <= 12'h72a; 
COS_ROM[3797] <= 12'h72b; 
COS_ROM[3798] <= 12'h72d; 
COS_ROM[3799] <= 12'h72e; 
COS_ROM[3800] <= 12'h730; 
COS_ROM[3801] <= 12'h731; 
COS_ROM[3802] <= 12'h732; 
COS_ROM[3803] <= 12'h734; 
COS_ROM[3804] <= 12'h735; 
COS_ROM[3805] <= 12'h736; 
COS_ROM[3806] <= 12'h738; 
COS_ROM[3807] <= 12'h739; 
COS_ROM[3808] <= 12'h73a; 
COS_ROM[3809] <= 12'h73c; 
COS_ROM[3810] <= 12'h73d; 
COS_ROM[3811] <= 12'h73e; 
COS_ROM[3812] <= 12'h740; 
COS_ROM[3813] <= 12'h741; 
COS_ROM[3814] <= 12'h742; 
COS_ROM[3815] <= 12'h744; 
COS_ROM[3816] <= 12'h745; 
COS_ROM[3817] <= 12'h746; 
COS_ROM[3818] <= 12'h748; 
COS_ROM[3819] <= 12'h749; 
COS_ROM[3820] <= 12'h74a; 
COS_ROM[3821] <= 12'h74c; 
COS_ROM[3822] <= 12'h74d; 
COS_ROM[3823] <= 12'h74e; 
COS_ROM[3824] <= 12'h74f; 
COS_ROM[3825] <= 12'h751; 
COS_ROM[3826] <= 12'h752; 
COS_ROM[3827] <= 12'h753; 
COS_ROM[3828] <= 12'h754; 
COS_ROM[3829] <= 12'h756; 
COS_ROM[3830] <= 12'h757; 
COS_ROM[3831] <= 12'h758; 
COS_ROM[3832] <= 12'h759; 
COS_ROM[3833] <= 12'h75b; 
COS_ROM[3834] <= 12'h75c; 
COS_ROM[3835] <= 12'h75d; 
COS_ROM[3836] <= 12'h75e; 
COS_ROM[3837] <= 12'h760; 
COS_ROM[3838] <= 12'h761; 
COS_ROM[3839] <= 12'h762; 
COS_ROM[3840] <= 12'h763; 
COS_ROM[3841] <= 12'h764; 
COS_ROM[3842] <= 12'h766; 
COS_ROM[3843] <= 12'h767; 
COS_ROM[3844] <= 12'h768; 
COS_ROM[3845] <= 12'h769; 
COS_ROM[3846] <= 12'h76a; 
COS_ROM[3847] <= 12'h76b; 
COS_ROM[3848] <= 12'h76d; 
COS_ROM[3849] <= 12'h76e; 
COS_ROM[3850] <= 12'h76f; 
COS_ROM[3851] <= 12'h770; 
COS_ROM[3852] <= 12'h771; 
COS_ROM[3853] <= 12'h772; 
COS_ROM[3854] <= 12'h774; 
COS_ROM[3855] <= 12'h775; 
COS_ROM[3856] <= 12'h776; 
COS_ROM[3857] <= 12'h777; 
COS_ROM[3858] <= 12'h778; 
COS_ROM[3859] <= 12'h779; 
COS_ROM[3860] <= 12'h77a; 
COS_ROM[3861] <= 12'h77b; 
COS_ROM[3862] <= 12'h77d; 
COS_ROM[3863] <= 12'h77e; 
COS_ROM[3864] <= 12'h77f; 
COS_ROM[3865] <= 12'h780; 
COS_ROM[3866] <= 12'h781; 
COS_ROM[3867] <= 12'h782; 
COS_ROM[3868] <= 12'h783; 
COS_ROM[3869] <= 12'h784; 
COS_ROM[3870] <= 12'h785; 
COS_ROM[3871] <= 12'h786; 
COS_ROM[3872] <= 12'h787; 
COS_ROM[3873] <= 12'h788; 
COS_ROM[3874] <= 12'h789; 
COS_ROM[3875] <= 12'h78a; 
COS_ROM[3876] <= 12'h78c; 
COS_ROM[3877] <= 12'h78d; 
COS_ROM[3878] <= 12'h78e; 
COS_ROM[3879] <= 12'h78f; 
COS_ROM[3880] <= 12'h790; 
COS_ROM[3881] <= 12'h791; 
COS_ROM[3882] <= 12'h792; 
COS_ROM[3883] <= 12'h793; 
COS_ROM[3884] <= 12'h794; 
COS_ROM[3885] <= 12'h795; 
COS_ROM[3886] <= 12'h796; 
COS_ROM[3887] <= 12'h797; 
COS_ROM[3888] <= 12'h798; 
COS_ROM[3889] <= 12'h799; 
COS_ROM[3890] <= 12'h79a; 
COS_ROM[3891] <= 12'h79b; 
COS_ROM[3892] <= 12'h79c; 
COS_ROM[3893] <= 12'h79d; 
COS_ROM[3894] <= 12'h79e; 
COS_ROM[3895] <= 12'h79e; 
COS_ROM[3896] <= 12'h79f; 
COS_ROM[3897] <= 12'h7a0; 
COS_ROM[3898] <= 12'h7a1; 
COS_ROM[3899] <= 12'h7a2; 
COS_ROM[3900] <= 12'h7a3; 
COS_ROM[3901] <= 12'h7a4; 
COS_ROM[3902] <= 12'h7a5; 
COS_ROM[3903] <= 12'h7a6; 
COS_ROM[3904] <= 12'h7a7; 
COS_ROM[3905] <= 12'h7a8; 
COS_ROM[3906] <= 12'h7a9; 
COS_ROM[3907] <= 12'h7aa; 
COS_ROM[3908] <= 12'h7aa; 
COS_ROM[3909] <= 12'h7ab; 
COS_ROM[3910] <= 12'h7ac; 
COS_ROM[3911] <= 12'h7ad; 
COS_ROM[3912] <= 12'h7ae; 
COS_ROM[3913] <= 12'h7af; 
COS_ROM[3914] <= 12'h7b0; 
COS_ROM[3915] <= 12'h7b1; 
COS_ROM[3916] <= 12'h7b1; 
COS_ROM[3917] <= 12'h7b2; 
COS_ROM[3918] <= 12'h7b3; 
COS_ROM[3919] <= 12'h7b4; 
COS_ROM[3920] <= 12'h7b5; 
COS_ROM[3921] <= 12'h7b6; 
COS_ROM[3922] <= 12'h7b7; 
COS_ROM[3923] <= 12'h7b7; 
COS_ROM[3924] <= 12'h7b8; 
COS_ROM[3925] <= 12'h7b9; 
COS_ROM[3926] <= 12'h7ba; 
COS_ROM[3927] <= 12'h7bb; 
COS_ROM[3928] <= 12'h7bb; 
COS_ROM[3929] <= 12'h7bc; 
COS_ROM[3930] <= 12'h7bd; 
COS_ROM[3931] <= 12'h7be; 
COS_ROM[3932] <= 12'h7bf; 
COS_ROM[3933] <= 12'h7bf; 
COS_ROM[3934] <= 12'h7c0; 
COS_ROM[3935] <= 12'h7c1; 
COS_ROM[3936] <= 12'h7c2; 
COS_ROM[3937] <= 12'h7c2; 
COS_ROM[3938] <= 12'h7c3; 
COS_ROM[3939] <= 12'h7c4; 
COS_ROM[3940] <= 12'h7c5; 
COS_ROM[3941] <= 12'h7c5; 
COS_ROM[3942] <= 12'h7c6; 
COS_ROM[3943] <= 12'h7c7; 
COS_ROM[3944] <= 12'h7c8; 
COS_ROM[3945] <= 12'h7c8; 
COS_ROM[3946] <= 12'h7c9; 
COS_ROM[3947] <= 12'h7ca; 
COS_ROM[3948] <= 12'h7ca; 
COS_ROM[3949] <= 12'h7cb; 
COS_ROM[3950] <= 12'h7cc; 
COS_ROM[3951] <= 12'h7cd; 
COS_ROM[3952] <= 12'h7cd; 
COS_ROM[3953] <= 12'h7ce; 
COS_ROM[3954] <= 12'h7cf; 
COS_ROM[3955] <= 12'h7cf; 
COS_ROM[3956] <= 12'h7d0; 
COS_ROM[3957] <= 12'h7d1; 
COS_ROM[3958] <= 12'h7d1; 
COS_ROM[3959] <= 12'h7d2; 
COS_ROM[3960] <= 12'h7d3; 
COS_ROM[3961] <= 12'h7d3; 
COS_ROM[3962] <= 12'h7d4; 
COS_ROM[3963] <= 12'h7d5; 
COS_ROM[3964] <= 12'h7d5; 
COS_ROM[3965] <= 12'h7d6; 
COS_ROM[3966] <= 12'h7d6; 
COS_ROM[3967] <= 12'h7d7; 
COS_ROM[3968] <= 12'h7d8; 
COS_ROM[3969] <= 12'h7d8; 
COS_ROM[3970] <= 12'h7d9; 
COS_ROM[3971] <= 12'h7d9; 
COS_ROM[3972] <= 12'h7da; 
COS_ROM[3973] <= 12'h7db; 
COS_ROM[3974] <= 12'h7db; 
COS_ROM[3975] <= 12'h7dc; 
COS_ROM[3976] <= 12'h7dc; 
COS_ROM[3977] <= 12'h7dd; 
COS_ROM[3978] <= 12'h7de; 
COS_ROM[3979] <= 12'h7de; 
COS_ROM[3980] <= 12'h7df; 
COS_ROM[3981] <= 12'h7df; 
COS_ROM[3982] <= 12'h7e0; 
COS_ROM[3983] <= 12'h7e0; 
COS_ROM[3984] <= 12'h7e1; 
COS_ROM[3985] <= 12'h7e1; 
COS_ROM[3986] <= 12'h7e2; 
COS_ROM[3987] <= 12'h7e2; 
COS_ROM[3988] <= 12'h7e3; 
COS_ROM[3989] <= 12'h7e3; 
COS_ROM[3990] <= 12'h7e4; 
COS_ROM[3991] <= 12'h7e5; 
COS_ROM[3992] <= 12'h7e5; 
COS_ROM[3993] <= 12'h7e6; 
COS_ROM[3994] <= 12'h7e6; 
COS_ROM[3995] <= 12'h7e6; 
COS_ROM[3996] <= 12'h7e7; 
COS_ROM[3997] <= 12'h7e7; 
COS_ROM[3998] <= 12'h7e8; 
COS_ROM[3999] <= 12'h7e8; 
COS_ROM[4000] <= 12'h7e9; 
COS_ROM[4001] <= 12'h7e9; 
COS_ROM[4002] <= 12'h7ea; 
COS_ROM[4003] <= 12'h7ea; 
COS_ROM[4004] <= 12'h7eb; 
COS_ROM[4005] <= 12'h7eb; 
COS_ROM[4006] <= 12'h7ec; 
COS_ROM[4007] <= 12'h7ec; 
COS_ROM[4008] <= 12'h7ec; 
COS_ROM[4009] <= 12'h7ed; 
COS_ROM[4010] <= 12'h7ed; 
COS_ROM[4011] <= 12'h7ee; 
COS_ROM[4012] <= 12'h7ee; 
COS_ROM[4013] <= 12'h7ee; 
COS_ROM[4014] <= 12'h7ef; 
COS_ROM[4015] <= 12'h7ef; 
COS_ROM[4016] <= 12'h7f0; 
COS_ROM[4017] <= 12'h7f0; 
COS_ROM[4018] <= 12'h7f0; 
COS_ROM[4019] <= 12'h7f1; 
COS_ROM[4020] <= 12'h7f1; 
COS_ROM[4021] <= 12'h7f1; 
COS_ROM[4022] <= 12'h7f2; 
COS_ROM[4023] <= 12'h7f2; 
COS_ROM[4024] <= 12'h7f3; 
COS_ROM[4025] <= 12'h7f3; 
COS_ROM[4026] <= 12'h7f3; 
COS_ROM[4027] <= 12'h7f4; 
COS_ROM[4028] <= 12'h7f4; 
COS_ROM[4029] <= 12'h7f4; 
COS_ROM[4030] <= 12'h7f5; 
COS_ROM[4031] <= 12'h7f5; 
COS_ROM[4032] <= 12'h7f5; 
COS_ROM[4033] <= 12'h7f5; 
COS_ROM[4034] <= 12'h7f6; 
COS_ROM[4035] <= 12'h7f6; 
COS_ROM[4036] <= 12'h7f6; 
COS_ROM[4037] <= 12'h7f7; 
COS_ROM[4038] <= 12'h7f7; 
COS_ROM[4039] <= 12'h7f7; 
COS_ROM[4040] <= 12'h7f7; 
COS_ROM[4041] <= 12'h7f8; 
COS_ROM[4042] <= 12'h7f8; 
COS_ROM[4043] <= 12'h7f8; 
COS_ROM[4044] <= 12'h7f8; 
COS_ROM[4045] <= 12'h7f9; 
COS_ROM[4046] <= 12'h7f9; 
COS_ROM[4047] <= 12'h7f9; 
COS_ROM[4048] <= 12'h7f9; 
COS_ROM[4049] <= 12'h7fa; 
COS_ROM[4050] <= 12'h7fa; 
COS_ROM[4051] <= 12'h7fa; 
COS_ROM[4052] <= 12'h7fa; 
COS_ROM[4053] <= 12'h7fb; 
COS_ROM[4054] <= 12'h7fb; 
COS_ROM[4055] <= 12'h7fb; 
COS_ROM[4056] <= 12'h7fb; 
COS_ROM[4057] <= 12'h7fb; 
COS_ROM[4058] <= 12'h7fc; 
COS_ROM[4059] <= 12'h7fc; 
COS_ROM[4060] <= 12'h7fc; 
COS_ROM[4061] <= 12'h7fc; 
COS_ROM[4062] <= 12'h7fc; 
COS_ROM[4063] <= 12'h7fc; 
COS_ROM[4064] <= 12'h7fd; 
COS_ROM[4065] <= 12'h7fd; 
COS_ROM[4066] <= 12'h7fd; 
COS_ROM[4067] <= 12'h7fd; 
COS_ROM[4068] <= 12'h7fd; 
COS_ROM[4069] <= 12'h7fd; 
COS_ROM[4070] <= 12'h7fd; 
COS_ROM[4071] <= 12'h7fd; 
COS_ROM[4072] <= 12'h7fe; 
COS_ROM[4073] <= 12'h7fe; 
COS_ROM[4074] <= 12'h7fe; 
COS_ROM[4075] <= 12'h7fe; 
COS_ROM[4076] <= 12'h7fe; 
COS_ROM[4077] <= 12'h7fe; 
COS_ROM[4078] <= 12'h7fe; 
COS_ROM[4079] <= 12'h7fe; 
COS_ROM[4080] <= 12'h7fe; 
COS_ROM[4081] <= 12'h7fe; 
COS_ROM[4082] <= 12'h7ff; 
COS_ROM[4083] <= 12'h7ff; 
COS_ROM[4084] <= 12'h7ff; 
COS_ROM[4085] <= 12'h7ff; 
COS_ROM[4086] <= 12'h7ff; 
COS_ROM[4087] <= 12'h7ff; 
COS_ROM[4088] <= 12'h7ff; 
COS_ROM[4089] <= 12'h7ff; 
COS_ROM[4090] <= 12'h7ff; 
COS_ROM[4091] <= 12'h7ff; 
COS_ROM[4092] <= 12'h7ff; 
COS_ROM[4093] <= 12'h7ff; 
COS_ROM[4094] <= 12'h7ff; 
COS_ROM[4095] <= 12'h7ff; 



end


endmodule

module waveform_gen (
    input wire clk,
	input wire reset,
    input wire en,
    input wire [31:0] phase_inc,
    output wire [11:0] sin_out,
    output wire [11:0] cos_out,
    output wire [11:0] squ_out,
	 output vco_out,
	 output desired_freq_sig);

// Phase accumulator and LUT address signals
reg [31:0] phase_acc;
wire [11:0] lut_addr;
reg [11:0] lut_addr_reg;
wire read;
// Sine/cosine LUT component instantiation
sincos_lut lut_inst (
    .clk(clk),
    .en(en),
    .addr(lut_addr),
    .sin_out(sin_out),
    .cos_out(cos_out)
);


// Phase accumulator logic
always @(posedge clk ) begin //or negedge reset
    if (~reset) begin
        phase_acc <= 32'b0;
    end else 
			if (en && ~read)
				begin
					phase_acc <= phase_acc + phase_inc;
				end
				else if(en&&read)
				begin
					phase_acc <= phase_acc + 32'h000D1B71;

				end
end

// Addressing the LUT using top 12 bits of the phase accumulator
assign lut_addr = phase_acc[31:20];
assign read = (phase_inc == 32'h000D1B71);


// Latency hiding registers for the LUT address
always @(posedge clk) begin

        lut_addr_reg <= lut_addr;

end

// Square wave output
assign squ_out = (lut_addr_reg[11]) ? 12'b011111111111 : 12'b100000000000;
assign vco_out = squ_out[11];

assign desired_freq_sig = read ? squ_out[11] : 1'b0;


endmodule
